// Generator : SpinalHDL dev    git head : 49a99dae7b6ed938ae50042417514f24dcaeaaa8
// Component : CoreNSCSCC
// Git hash  : 63ae007975c3d36491b8fbaf9c85d0550b9457d0

`timescale 1ns/1ps

module CoreNSCSCC (
  input  wire          clk,
  output wire [7:0]    io_dpy0,
  output wire [7:0]    io_dpy1,
  output wire [15:0]   io_leds,
  input  wire          io_switch_btn,
  input  wire [31:0]   io_isram_dout,
  output wire [19:0]   io_isram_addr,
  output wire [31:0]   io_isram_din,
  output wire          io_isram_en,
  output wire          io_isram_re,
  output wire          io_isram_we,
  output wire [3:0]    io_isram_wmask,
  input  wire [31:0]   io_dsram_dout,
  output wire [19:0]   io_dsram_addr,
  output wire [31:0]   io_dsram_din,
  output wire          io_dsram_en,
  output wire          io_dsram_re,
  output wire          io_dsram_we,
  output wire [3:0]    io_dsram_wmask,
  input  wire          io_uart_ar_ready,
  input  wire [7:0]    io_uart_r_bits_id,
  input  wire [1:0]    io_uart_r_bits_resp,
  input  wire [31:0]   io_uart_r_bits_data,
  input  wire          io_uart_r_bits_last,
  input  wire          io_uart_r_valid,
  input  wire          io_uart_aw_ready,
  input  wire          io_uart_w_ready,
  input  wire [7:0]    io_uart_b_bits_id,
  input  wire [1:0]    io_uart_b_bits_resp,
  input  wire          io_uart_b_valid,
  output wire [7:0]    io_uart_ar_bits_id,
  output wire [31:0]   io_uart_ar_bits_addr,
  output wire [7:0]    io_uart_ar_bits_len,
  output wire [2:0]    io_uart_ar_bits_size,
  output wire [1:0]    io_uart_ar_bits_burst,
  output wire          io_uart_ar_valid,
  output wire          io_uart_r_ready,
  output wire [7:0]    io_uart_aw_bits_id,
  output wire [31:0]   io_uart_aw_bits_addr,
  output wire [7:0]    io_uart_aw_bits_len,
  output wire [2:0]    io_uart_aw_bits_size,
  output wire [1:0]    io_uart_aw_bits_burst,
  output wire          io_uart_aw_valid,
  output wire [31:0]   io_uart_w_bits_data,
  output wire [3:0]    io_uart_w_bits_strb,
  output wire          io_uart_w_bits_last,
  output wire          io_uart_w_valid,
  output wire          io_uart_b_ready,
  input  wire          reset
);
  localparam BranchCondition_NUL = 5'd0;
  localparam BranchCondition_EQ = 5'd1;
  localparam BranchCondition_NE = 5'd2;
  localparam BranchCondition_LT = 5'd3;
  localparam BranchCondition_GE = 5'd4;
  localparam BranchCondition_LTU = 5'd5;
  localparam BranchCondition_GEU = 5'd6;
  localparam BranchCondition_EQZ = 5'd7;
  localparam BranchCondition_NEZ = 5'd8;
  localparam BranchCondition_LTZ = 5'd9;
  localparam BranchCondition_GEZ = 5'd10;
  localparam BranchCondition_GTZ = 5'd11;
  localparam BranchCondition_LEZ = 5'd12;
  localparam BranchCondition_F_EQ = 5'd13;
  localparam BranchCondition_F_NE = 5'd14;
  localparam BranchCondition_F_LT = 5'd15;
  localparam BranchCondition_F_LE = 5'd16;
  localparam BranchCondition_F_UN = 5'd17;
  localparam BranchCondition_LA_CF_TRUE = 5'd18;
  localparam BranchCondition_LA_CF_FALSE = 5'd19;
  localparam ArchRegType_GPR = 2'd0;
  localparam ArchRegType_FPR = 2'd1;
  localparam ArchRegType_CSR = 2'd2;
  localparam ArchRegType_LA_CF = 2'd3;
  localparam IntAluExceptionCode_NONE = 1'd0;
  localparam IntAluExceptionCode_UNDEFINED_ALU_OP = 1'd1;
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam BaseUopCode_NOP = 5'd0;
  localparam BaseUopCode_ILLEGAL = 5'd1;
  localparam BaseUopCode_ALU = 5'd2;
  localparam BaseUopCode_SHIFT = 5'd3;
  localparam BaseUopCode_MUL = 5'd4;
  localparam BaseUopCode_DIV = 5'd5;
  localparam BaseUopCode_LOAD = 5'd6;
  localparam BaseUopCode_STORE = 5'd7;
  localparam BaseUopCode_ATOMIC = 5'd8;
  localparam BaseUopCode_MEM_BARRIER = 5'd9;
  localparam BaseUopCode_PREFETCH = 5'd10;
  localparam BaseUopCode_BRANCH = 5'd11;
  localparam BaseUopCode_JUMP_REG = 5'd12;
  localparam BaseUopCode_JUMP_IMM = 5'd13;
  localparam BaseUopCode_SYSTEM_OP = 5'd14;
  localparam BaseUopCode_CSR_ACCESS = 5'd15;
  localparam BaseUopCode_FPU_ALU = 5'd16;
  localparam BaseUopCode_FPU_CVT = 5'd17;
  localparam BaseUopCode_FPU_CMP = 5'd18;
  localparam BaseUopCode_FPU_SEL = 5'd19;
  localparam BaseUopCode_LA_BITMANIP = 5'd20;
  localparam BaseUopCode_LA_CACOP = 5'd21;
  localparam BaseUopCode_LA_TLB = 5'd22;
  localparam BaseUopCode_IDLE = 5'd23;
  localparam ExeUnitType_NONE = 4'd0;
  localparam ExeUnitType_ALU_INT = 4'd1;
  localparam ExeUnitType_MUL_INT = 4'd2;
  localparam ExeUnitType_DIV_INT = 4'd3;
  localparam ExeUnitType_MEM = 4'd4;
  localparam ExeUnitType_BRU = 4'd5;
  localparam ExeUnitType_CSR = 4'd6;
  localparam ExeUnitType_FPU_ADD_MUL_CVT_CMP = 4'd7;
  localparam ExeUnitType_FPU_DIV_SQRT = 4'd8;
  localparam IsaType_UNKNOWN = 2'd0;
  localparam IsaType_DEMO = 2'd1;
  localparam IsaType_RISCV = 2'd2;
  localparam IsaType_LOONGARCH = 2'd3;
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;
  localparam DecodeExCode_INVALID = 2'd0;
  localparam DecodeExCode_FETCH_ERROR = 2'd1;
  localparam DecodeExCode_DECODE_ERROR = 2'd2;
  localparam DecodeExCode_OK = 2'd3;
  localparam FlushReason_NONE = 2'd0;
  localparam FlushReason_FULL_FLUSH = 2'd1;
  localparam FlushReason_ROLLBACK_TO_ROB_IDX = 2'd2;
  localparam ICachePlugin_logic_refill_fsm_BOOT = 5'd1;
  localparam ICachePlugin_logic_refill_fsm_IDLE = 5'd2;
  localparam ICachePlugin_logic_refill_fsm_SEND_REQ = 5'd4;
  localparam ICachePlugin_logic_refill_fsm_RECEIVE_DATA = 5'd8;
  localparam ICachePlugin_logic_refill_fsm_COMMIT = 5'd16;
  localparam ICachePlugin_logic_refill_fsm_BOOT_OH_ID = 0;
  localparam ICachePlugin_logic_refill_fsm_IDLE_OH_ID = 1;
  localparam ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID = 2;
  localparam ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID = 3;
  localparam ICachePlugin_logic_refill_fsm_COMMIT_OH_ID = 4;

  reg                 DataCachePlugin_setup_cache_io_mem_read_cmd_ready;
  wire                DataCachePlugin_setup_cache_io_mem_read_rsp_payload_error;
  reg                 DataCachePlugin_setup_cache_io_mem_write_cmd_ready;
  wire                DataCachePlugin_setup_cache_io_mem_write_rsp_payload_error;
  wire                oneShot_13_io_triggerIn;
  wire                ROBPlugin_robComponent_io_allocate_0_valid;
  reg                 ROBPlugin_robComponent_io_writeback_4_fire;
  reg        [3:0]    ROBPlugin_robComponent_io_writeback_4_robPtr;
  reg        [31:0]   ROBPlugin_robComponent_io_writeback_4_result;
  reg                 ROBPlugin_robComponent_io_writeback_4_exceptionOccurred;
  reg        [7:0]    ROBPlugin_robComponent_io_writeback_4_exceptionCodeIn;
  wire                RenameMapTablePlugin_early_setup_rat_io_writePorts_0_wen;
  reg                 RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_valid;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_0;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_1;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_2;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_3;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_4;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_5;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_6;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_7;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_8;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_9;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_10;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_11;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_12;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_13;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_14;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_15;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_16;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_17;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_18;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_19;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_20;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_21;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_22;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_23;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_24;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_25;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_26;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_27;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_28;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_29;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_30;
  reg        [5:0]    RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_31;
  wire                SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_enable;
  reg                 SimpleFreeListPlugin_early_setup_freeList_io_recover;
  wire                oneShot_14_io_triggerIn;
  wire                oneShot_15_io_triggerIn;
  wire                oneShot_16_io_triggerIn;
  wire                oneShot_17_io_triggerIn;
  wire                DebugDisplayPlugin_hw_dpyController_io_dp0;
  wire                oneShot_18_io_triggerIn;
  wire       [31:0]   lA32RSimpleDecoder_1_io_pcIn;
  wire                oneShot_20_io_triggerIn;
  wire                oneShot_21_io_triggerIn;
  wire       [31:0]   multiplierBlackbox_A;
  wire       [31:0]   multiplierBlackbox_B;
  wire                oneShot_22_io_triggerIn;
  wire                oneShot_23_io_triggerIn;
  wire       [0:0]    streamDemux_1_io_select;
  wire                oneShot_24_io_triggerIn;
  wire                oneShot_25_io_triggerIn;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_valid;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_pc;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_0;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_1;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_2;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_3;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isBranch;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isJump;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isDirectJump;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_jumpOffset;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isIdle;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isBranch;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isJump;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isDirectJump;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_jumpOffset;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isIdle;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isBranch;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isJump;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isDirectJump;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_jumpOffset;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isIdle;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isBranch;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isJump;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isDirectJump;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_jumpOffset;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isIdle;
  reg        [3:0]    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_branchMask;
  reg                 FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_fault;
  reg        [2:0]    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_numValidInstructions;
  reg        [1:0]    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_startInstructionIndex;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_ready;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_flush;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_instruction;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_instruction;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_instruction;
  reg        [31:0]   FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_instruction;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_ready;
  wire       [3:0]    io_axiOut_readOnly_decoder_io_outputs_0_r_payload_id;
  wire       [3:0]    io_axiOut_readOnly_decoder_io_outputs_1_r_payload_id;
  wire       [3:0]    io_axiOut_readOnly_decoder_io_outputs_2_r_payload_id;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_0_b_payload_id;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_1_b_payload_id;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_2_b_payload_id;
  wire       [3:0]    io_axiOut_readOnly_decoder_1_io_outputs_0_r_payload_id;
  wire       [3:0]    io_axiOut_readOnly_decoder_1_io_outputs_1_r_payload_id;
  wire       [3:0]    io_axiOut_readOnly_decoder_1_io_outputs_2_r_payload_id;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_0_b_payload_id;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_1_b_payload_id;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_2_b_payload_id;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_r_payload_id;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_r_payload_id;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_r_payload_id;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_b_payload_id;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_b_payload_id;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_b_payload_id;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_r_payload_id;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_r_payload_id;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_r_payload_id;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_b_payload_id;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_b_payload_id;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_b_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_3_io_inputs_0_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_3_io_inputs_1_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_3_io_inputs_2_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_3_io_inputs_3_ar_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_3_io_inputs_0_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_3_io_inputs_1_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_3_io_inputs_2_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_3_io_inputs_3_aw_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_4_io_inputs_0_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_4_io_inputs_1_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_4_io_inputs_2_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_4_io_inputs_3_ar_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_4_io_inputs_0_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_4_io_inputs_1_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_4_io_inputs_2_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_4_io_inputs_3_aw_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_5_io_inputs_0_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_5_io_inputs_1_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_5_io_inputs_2_ar_payload_id;
  wire       [4:0]    axi4ReadOnlyArbiter_5_io_inputs_3_ar_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_5_io_inputs_0_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_5_io_inputs_1_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_5_io_inputs_2_aw_payload_id;
  wire       [4:0]    axi4WriteOnlyArbiter_5_io_inputs_3_aw_payload_id;
  reg        [42:0]   ICachePlugin_logic_storage_tagLruRam_spinal_port1;
  reg        [127:0]  ICachePlugin_logic_storage_dataRams_0_spinal_port0;
  reg        [127:0]  ICachePlugin_logic_storage_dataRams_1_spinal_port0;
  reg        [1:0]    BpuPipelinePlugin_logic_pht_spinal_port0;
  reg        [1:0]    BpuPipelinePlugin_logic_pht_spinal_port1;
  reg        [54:0]   BpuPipelinePlugin_logic_btb_spinal_port0;
  wire                AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_valid;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_data;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_physDest_idx;
  wire                AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_writesToPhysReg;
  wire       [3:0]    AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_robPtr;
  wire                AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_hasException;
  wire       [0:0]    AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_exceptionCode;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_axi_ar_ready;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_axi_aw_ready;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_axi_w_ready;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_valid;
  wire       [31:0]   CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_data;
  wire       [6:0]    CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_id;
  wire       [1:0]    CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_resp;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_last;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_valid;
  wire       [6:0]    CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_payload_id;
  wire       [1:0]    CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_payload_resp;
  wire       [31:0]   CoreMemSysPlugin_hw_baseramCtrl_io_ram_data_write;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_ram_data_writeEnable;
  wire       [19:0]   CoreMemSysPlugin_hw_baseramCtrl_io_ram_addr;
  wire       [3:0]    CoreMemSysPlugin_hw_baseramCtrl_io_ram_be_n;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_ram_ce_n;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_ram_oe_n;
  wire                CoreMemSysPlugin_hw_baseramCtrl_io_ram_we_n;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_axi_ar_ready;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_axi_aw_ready;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_axi_w_ready;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_axi_r_valid;
  wire       [31:0]   CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_data;
  wire       [6:0]    CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_id;
  wire       [1:0]    CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_resp;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_last;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_axi_b_valid;
  wire       [6:0]    CoreMemSysPlugin_hw_extramCtrl_io_axi_b_payload_id;
  wire       [1:0]    CoreMemSysPlugin_hw_extramCtrl_io_axi_b_payload_resp;
  wire       [31:0]   CoreMemSysPlugin_hw_extramCtrl_io_ram_data_write;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_ram_data_writeEnable;
  wire       [19:0]   CoreMemSysPlugin_hw_extramCtrl_io_ram_addr;
  wire       [3:0]    CoreMemSysPlugin_hw_extramCtrl_io_ram_be_n;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_ram_ce_n;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_ram_oe_n;
  wire                CoreMemSysPlugin_hw_extramCtrl_io_ram_we_n;
  wire                DataCachePlugin_setup_cache_io_load_cmd_ready;
  wire                DataCachePlugin_setup_cache_io_load_rsp_valid;
  wire       [31:0]   DataCachePlugin_setup_cache_io_load_rsp_payload_data;
  wire                DataCachePlugin_setup_cache_io_load_rsp_payload_fault;
  wire                DataCachePlugin_setup_cache_io_load_rsp_payload_redo;
  wire       [7:0]    DataCachePlugin_setup_cache_io_load_rsp_payload_refillSlot;
  wire                DataCachePlugin_setup_cache_io_load_rsp_payload_refillSlotAny;
  wire       [2:0]    DataCachePlugin_setup_cache_io_load_rsp_payload_id;
  wire                DataCachePlugin_setup_cache_io_store_cmd_ready;
  wire                DataCachePlugin_setup_cache_io_store_rsp_valid;
  wire                DataCachePlugin_setup_cache_io_store_rsp_payload_fault;
  wire                DataCachePlugin_setup_cache_io_store_rsp_payload_redo;
  wire       [7:0]    DataCachePlugin_setup_cache_io_store_rsp_payload_refillSlot;
  wire                DataCachePlugin_setup_cache_io_store_rsp_payload_refillSlotAny;
  wire                DataCachePlugin_setup_cache_io_store_rsp_payload_flush;
  wire                DataCachePlugin_setup_cache_io_store_rsp_payload_prefetch;
  wire       [31:0]   DataCachePlugin_setup_cache_io_store_rsp_payload_address;
  wire                DataCachePlugin_setup_cache_io_store_rsp_payload_io;
  wire       [2:0]    DataCachePlugin_setup_cache_io_store_rsp_payload_id;
  wire                DataCachePlugin_setup_cache_io_mem_read_cmd_valid;
  wire       [2:0]    DataCachePlugin_setup_cache_io_mem_read_cmd_payload_id;
  wire       [31:0]   DataCachePlugin_setup_cache_io_mem_read_cmd_payload_address;
  wire                DataCachePlugin_setup_cache_io_mem_read_rsp_ready;
  wire                DataCachePlugin_setup_cache_io_mem_write_cmd_valid;
  wire                DataCachePlugin_setup_cache_io_mem_write_cmd_payload_last;
  wire       [31:0]   DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_address;
  wire       [31:0]   DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_data;
  wire       [2:0]    DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_id;
  wire       [7:0]    DataCachePlugin_setup_cache_io_refillCompletions;
  wire                DataCachePlugin_setup_cache_io_refillEvent;
  wire                DataCachePlugin_setup_cache_io_writebackEvent;
  wire                DataCachePlugin_setup_cache_io_writebackBusy;
  wire                oneShot_13_io_pulseOut;
  wire                FetchPipelinePlugin_setup_fetchOutput_io_push_ready;
  wire                FetchPipelinePlugin_setup_fetchOutput_io_pop_valid;
  wire       [31:0]   FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_pc;
  wire       [31:0]   FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_instruction;
  wire                FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_isBranch;
  wire                FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_isJump;
  wire                FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_jumpOffset;
  wire                FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_isIdle;
  wire                FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_isTaken;
  wire       [31:0]   FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_target;
  wire                FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_wasPredicted;
  wire       [2:0]    FetchPipelinePlugin_setup_fetchOutput_io_occupancy;
  wire       [2:0]    FetchPipelinePlugin_setup_fetchOutput_io_availability;
  wire       [3:0]    ROBPlugin_robComponent_io_allocate_0_robPtr;
  wire                ROBPlugin_robComponent_io_allocate_0_ready;
  wire                ROBPlugin_robComponent_io_canAllocate_0;
  wire                ROBPlugin_robComponent_io_commit_0_valid;
  wire                ROBPlugin_robComponent_io_commit_0_canCommit;
  wire       [31:0]   ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_pc;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isValid;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_uopCode;
  wire       [3:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_exeUnit;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isa;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archDest_idx;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archDest_rtype;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_writeArchDestEn;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archSrc1_idx;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_useArchSrc1;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archSrc2_idx;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_useArchSrc2;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_usePcForAddr;
  wire       [31:0]   ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_imm;
  wire       [2:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_immUsage;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_isSub;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_isAdd;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_isSigned;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRight;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_isArithmetic;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRotate;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_isDoubleWord;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isDiv;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isSigned;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isWordOp;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_size;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isStore;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isLoadLinked;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isStoreCond;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_atomicOp;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isFence;
  wire       [7:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_fenceMode;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isCacheOp;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_cacheOpType;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isPrefetch;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_isLink;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_isIndirect;
  wire       [2:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_laCfIdx;
  wire       [3:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest;
  wire       [2:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_roundingMode;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_isIntegerDest;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_isSignedCvt;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fcmpCond;
  wire       [13:0]   ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_isWrite;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_isRead;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_isExchange;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  wire       [19:0]   ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_sysCtrl_isExceptionReturn;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_sysCtrl_isTlbOp;
  wire       [3:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_sysCtrl_tlbOpType;
  wire       [1:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_hasDecodeException;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isMicrocode;
  wire       [7:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_microcodeEntry;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isSerializing;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isBranchOrJump;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken;
  wire       [31:0]   ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchPrediction_target;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchPrediction_wasPredicted;
  wire       [5:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physSrc1_idx;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physSrc1IsFpr;
  wire       [5:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physSrc2_idx;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physSrc2IsFpr;
  wire       [5:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physDest_idx;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physDestIsFpr;
  wire       [5:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_oldPhysDest_idx;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_oldPhysDestIsFpr;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_allocatesPhysDest;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_writesToPhysReg;
  wire       [3:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_robPtr;
  wire       [15:0]   ROBPlugin_robComponent_io_commit_0_entry_payload_uop_uniqueId;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_dispatched;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_executed;
  wire                ROBPlugin_robComponent_io_commit_0_entry_payload_uop_hasException;
  wire       [7:0]    ROBPlugin_robComponent_io_commit_0_entry_payload_uop_exceptionCode;
  wire       [31:0]   ROBPlugin_robComponent_io_commit_0_entry_payload_pc;
  wire                ROBPlugin_robComponent_io_commit_0_entry_status_busy;
  wire                ROBPlugin_robComponent_io_commit_0_entry_status_done;
  wire                ROBPlugin_robComponent_io_commit_0_entry_status_isMispredictedBranch;
  wire                ROBPlugin_robComponent_io_commit_0_entry_status_isTaken;
  wire       [31:0]   ROBPlugin_robComponent_io_commit_0_entry_status_result;
  wire                ROBPlugin_robComponent_io_commit_0_entry_status_hasException;
  wire       [7:0]    ROBPlugin_robComponent_io_commit_0_entry_status_exceptionCode;
  wire                ROBPlugin_robComponent_io_commit_0_entry_status_genBit;
  wire                ROBPlugin_robComponent_io_flushed;
  wire                ROBPlugin_robComponent_io_empty;
  wire       [3:0]    ROBPlugin_robComponent_io_headPtrOut;
  wire       [3:0]    ROBPlugin_robComponent_io_tailPtrOut;
  wire       [3:0]    ROBPlugin_robComponent_io_countOut;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_readPorts_0_physReg;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_readPorts_1_physReg;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_readPorts_2_physReg;
  wire                RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_ready;
  wire                RenameMapTablePlugin_early_setup_rat_io_checkpointSave_ready;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_0;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_1;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_2;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_3;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_4;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_5;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_6;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_7;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_8;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_9;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_10;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_11;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_12;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_13;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_14;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_15;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_16;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_17;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_18;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_19;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_20;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_21;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_22;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_23;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_24;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_25;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_26;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_27;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_28;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_29;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_30;
  wire       [5:0]    RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_31;
  wire       [5:0]    SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_physReg;
  wire                SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_success;
  wire       [5:0]    SimpleFreeListPlugin_early_setup_freeList_io_numFreeRegs;
  wire                oneShot_14_io_pulseOut;
  wire                oneShot_15_io_pulseOut;
  wire                oneShot_16_io_pulseOut;
  wire                oneShot_17_io_pulseOut;
  wire       [31:0]   RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_pc;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isValid;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_uopCode;
  wire       [3:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_exeUnit;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isa;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archDest_idx;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archDest_rtype;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_writeArchDestEn;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc1_idx;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc1_rtype;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_useArchSrc1;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc2_idx;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc2_rtype;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_useArchSrc2;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_usePcForAddr;
  wire       [31:0]   RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_imm;
  wire       [2:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_immUsage;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_valid;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isSub;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isAdd;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isSigned;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_logicOp;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_valid;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isRight;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isArithmetic;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isRotate;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isDoubleWord;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_valid;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isDiv;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isSigned;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isWordOp;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_size;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isSignedLoad;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isStore;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isLoadLinked;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isStoreCond;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_atomicOp;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isFence;
  wire       [7:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_fenceMode;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isCacheOp;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_cacheOpType;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isPrefetch;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_condition;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isJump;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isLink;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isIndirect;
  wire       [2:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_laCfIdx;
  wire       [3:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_opType;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest;
  wire       [2:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_roundingMode;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_isIntegerDest;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_isSignedCvt;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fcmpCond;
  wire       [13:0]   RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_csrAddr;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isWrite;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isRead;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isExchange;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_useUimmAsSrc;
  wire       [19:0]   RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_sysCode;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_isExceptionReturn;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_isTlbOp;
  wire       [3:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_tlbOpType;
  wire       [1:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_decodeExceptionCode;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_hasDecodeException;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isMicrocode;
  wire       [7:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_microcodeEntry;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isSerializing;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isBranchOrJump;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_isTaken;
  wire       [31:0]   RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_target;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_wasPredicted;
  wire       [5:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc1_idx;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc1IsFpr;
  wire       [5:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc2_idx;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc2IsFpr;
  wire       [5:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physDest_idx;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physDestIsFpr;
  wire       [5:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_oldPhysDest_idx;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_oldPhysDestIsFpr;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_allocatesPhysDest;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_writesToPhysReg;
  wire       [3:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_robPtr;
  wire       [15:0]   RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_uniqueId;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_dispatched;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_executed;
  wire                RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_hasException;
  wire       [7:0]    RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_exceptionCode;
  wire       [0:0]    RenamePlugin_setup_renameUnit_io_numPhysRegsRequired;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_ratReadPorts_0_archReg;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_ratReadPorts_1_archReg;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_ratReadPorts_2_archReg;
  wire                RenamePlugin_setup_renameUnit_io_ratWritePorts_0_wen;
  wire       [4:0]    RenamePlugin_setup_renameUnit_io_ratWritePorts_0_archReg;
  wire       [5:0]    RenamePlugin_setup_renameUnit_io_ratWritePorts_0_physReg;
  wire       [7:0]    DebugDisplayPlugin_hw_dpyController_io_dpy0_out;
  wire       [7:0]    DebugDisplayPlugin_hw_dpyController_io_dpy1_out;
  wire                streamArbiter_8_io_inputs_0_ready;
  wire                streamArbiter_8_io_inputs_1_ready;
  wire                streamArbiter_8_io_inputs_2_ready;
  wire                streamArbiter_8_io_output_valid;
  wire       [5:0]    streamArbiter_8_io_output_payload_physRegIdx;
  wire       [31:0]   streamArbiter_8_io_output_payload_physRegData;
  wire       [3:0]    streamArbiter_8_io_output_payload_robPtr;
  wire                streamArbiter_8_io_output_payload_isFPR;
  wire                streamArbiter_8_io_output_payload_hasException;
  wire       [7:0]    streamArbiter_8_io_output_payload_exceptionCode;
  wire       [1:0]    streamArbiter_8_io_chosen;
  wire       [2:0]    streamArbiter_8_io_chosenOH;
  wire                oneShot_18_io_pulseOut;
  wire                oneShot_19_io_pulseOut;
  wire       [31:0]   lA32RSimpleDecoder_1_io_decodedUop_pc;
  wire                lA32RSimpleDecoder_1_io_decodedUop_isValid;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_uopCode;
  wire       [3:0]    lA32RSimpleDecoder_1_io_decodedUop_exeUnit;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_isa;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_archDest_idx;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_archDest_rtype;
  wire                lA32RSimpleDecoder_1_io_decodedUop_writeArchDestEn;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_archSrc1_idx;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_archSrc1_rtype;
  wire                lA32RSimpleDecoder_1_io_decodedUop_useArchSrc1;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_archSrc2_idx;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_archSrc2_rtype;
  wire                lA32RSimpleDecoder_1_io_decodedUop_useArchSrc2;
  wire                lA32RSimpleDecoder_1_io_decodedUop_usePcForAddr;
  wire       [31:0]   lA32RSimpleDecoder_1_io_decodedUop_imm;
  wire       [2:0]    lA32RSimpleDecoder_1_io_decodedUop_immUsage;
  wire                lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_valid;
  wire                lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isSub;
  wire                lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isAdd;
  wire                lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isSigned;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_logicOp;
  wire                lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_valid;
  wire                lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isRight;
  wire                lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isArithmetic;
  wire                lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isRotate;
  wire                lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isDoubleWord;
  wire                lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_valid;
  wire                lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isDiv;
  wire                lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isSigned;
  wire                lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isWordOp;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_memCtrl_size;
  wire                lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isSignedLoad;
  wire                lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isStore;
  wire                lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isLoadLinked;
  wire                lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isStoreCond;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_memCtrl_atomicOp;
  wire                lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isFence;
  wire       [7:0]    lA32RSimpleDecoder_1_io_decodedUop_memCtrl_fenceMode;
  wire                lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isCacheOp;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_memCtrl_cacheOpType;
  wire                lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isPrefetch;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_condition;
  wire                lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isJump;
  wire                lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isLink;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_linkReg_idx;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_linkReg_rtype;
  wire                lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isIndirect;
  wire       [2:0]    lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_laCfIdx;
  wire       [3:0]    lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_opType;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeDest;
  wire       [2:0]    lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_roundingMode;
  wire                lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_isIntegerDest;
  wire                lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_isSignedCvt;
  wire                lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fcmpCond;
  wire       [13:0]   lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_csrAddr;
  wire                lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isWrite;
  wire                lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isRead;
  wire                lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isExchange;
  wire                lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_useUimmAsSrc;
  wire       [19:0]   lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_sysCode;
  wire                lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_isExceptionReturn;
  wire                lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_isTlbOp;
  wire       [3:0]    lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_tlbOpType;
  wire       [1:0]    lA32RSimpleDecoder_1_io_decodedUop_decodeExceptionCode;
  wire                lA32RSimpleDecoder_1_io_decodedUop_hasDecodeException;
  wire                lA32RSimpleDecoder_1_io_decodedUop_isMicrocode;
  wire       [7:0]    lA32RSimpleDecoder_1_io_decodedUop_microcodeEntry;
  wire                lA32RSimpleDecoder_1_io_decodedUop_isSerializing;
  wire                lA32RSimpleDecoder_1_io_decodedUop_isBranchOrJump;
  wire                lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_isTaken;
  wire       [31:0]   lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_target;
  wire                lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_wasPredicted;
  wire                issueQueueComponent_4_io_allocateIn_ready;
  wire                issueQueueComponent_4_io_issueOut_valid;
  wire       [3:0]    issueQueueComponent_4_io_issueOut_payload_robPtr;
  wire       [5:0]    issueQueueComponent_4_io_issueOut_payload_physDest_idx;
  wire                issueQueueComponent_4_io_issueOut_payload_physDestIsFpr;
  wire                issueQueueComponent_4_io_issueOut_payload_writesToPhysReg;
  wire                issueQueueComponent_4_io_issueOut_payload_useSrc1;
  wire       [31:0]   issueQueueComponent_4_io_issueOut_payload_src1Data;
  wire       [5:0]    issueQueueComponent_4_io_issueOut_payload_src1Tag;
  wire                issueQueueComponent_4_io_issueOut_payload_src1Ready;
  wire                issueQueueComponent_4_io_issueOut_payload_src1IsFpr;
  wire                issueQueueComponent_4_io_issueOut_payload_useSrc2;
  wire       [31:0]   issueQueueComponent_4_io_issueOut_payload_src2Data;
  wire       [5:0]    issueQueueComponent_4_io_issueOut_payload_src2Tag;
  wire                issueQueueComponent_4_io_issueOut_payload_src2Ready;
  wire                issueQueueComponent_4_io_issueOut_payload_src2IsFpr;
  wire                issueQueueComponent_4_io_issueOut_payload_aluCtrl_valid;
  wire                issueQueueComponent_4_io_issueOut_payload_aluCtrl_isSub;
  wire                issueQueueComponent_4_io_issueOut_payload_aluCtrl_isAdd;
  wire                issueQueueComponent_4_io_issueOut_payload_aluCtrl_isSigned;
  wire       [1:0]    issueQueueComponent_4_io_issueOut_payload_aluCtrl_logicOp;
  wire                issueQueueComponent_4_io_issueOut_payload_shiftCtrl_valid;
  wire                issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isRight;
  wire                issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isArithmetic;
  wire                issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isRotate;
  wire                issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isDoubleWord;
  wire       [31:0]   issueQueueComponent_4_io_issueOut_payload_imm;
  wire       [2:0]    issueQueueComponent_4_io_issueOut_payload_immUsage;
  wire                issueQueueComponent_5_io_allocateIn_ready;
  wire                issueQueueComponent_5_io_issueOut_valid;
  wire       [31:0]   issueQueueComponent_5_io_issueOut_payload_uop_decoded_pc;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_isValid;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_uopCode;
  wire       [3:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_exeUnit;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_isa;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_archDest_idx;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_archDest_rtype;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_writeArchDestEn;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc1_idx;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc1_rtype;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_useArchSrc1;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc2_idx;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc2_rtype;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_useArchSrc2;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_usePcForAddr;
  wire       [31:0]   issueQueueComponent_5_io_issueOut_payload_uop_decoded_imm;
  wire       [2:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_immUsage;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_valid;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isSub;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isAdd;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isSigned;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_logicOp;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_valid;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isRight;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_valid;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_size;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isStore;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_atomicOp;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isFence;
  wire       [7:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_fenceMode;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_condition;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isJump;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isLink;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect;
  wire       [2:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx;
  wire       [3:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_opType;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest;
  wire       [2:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond;
  wire       [13:0]   issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isWrite;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isRead;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isExchange;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  wire       [19:0]   issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_sysCode;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp;
  wire       [3:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType;
  wire       [1:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_decodeExceptionCode;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_hasDecodeException;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_isMicrocode;
  wire       [7:0]    issueQueueComponent_5_io_issueOut_payload_uop_decoded_microcodeEntry;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_isSerializing;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_isBranchOrJump;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_isTaken;
  wire       [31:0]   issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_target;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted;
  wire       [5:0]    issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc1_idx;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc1IsFpr;
  wire       [5:0]    issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc2_idx;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc2IsFpr;
  wire       [5:0]    issueQueueComponent_5_io_issueOut_payload_uop_rename_physDest_idx;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_rename_physDestIsFpr;
  wire       [5:0]    issueQueueComponent_5_io_issueOut_payload_uop_rename_oldPhysDest_idx;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_rename_oldPhysDestIsFpr;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_rename_allocatesPhysDest;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_rename_writesToPhysReg;
  wire       [3:0]    issueQueueComponent_5_io_issueOut_payload_uop_robPtr;
  wire       [15:0]   issueQueueComponent_5_io_issueOut_payload_uop_uniqueId;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_dispatched;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_executed;
  wire                issueQueueComponent_5_io_issueOut_payload_uop_hasException;
  wire       [7:0]    issueQueueComponent_5_io_issueOut_payload_uop_exceptionCode;
  wire       [3:0]    issueQueueComponent_5_io_issueOut_payload_robPtr;
  wire       [5:0]    issueQueueComponent_5_io_issueOut_payload_physDest_idx;
  wire                issueQueueComponent_5_io_issueOut_payload_physDestIsFpr;
  wire                issueQueueComponent_5_io_issueOut_payload_writesToPhysReg;
  wire                issueQueueComponent_5_io_issueOut_payload_useSrc1;
  wire       [31:0]   issueQueueComponent_5_io_issueOut_payload_src1Data;
  wire       [5:0]    issueQueueComponent_5_io_issueOut_payload_src1Tag;
  wire                issueQueueComponent_5_io_issueOut_payload_src1Ready;
  wire                issueQueueComponent_5_io_issueOut_payload_src1IsFpr;
  wire                issueQueueComponent_5_io_issueOut_payload_useSrc2;
  wire       [31:0]   issueQueueComponent_5_io_issueOut_payload_src2Data;
  wire       [5:0]    issueQueueComponent_5_io_issueOut_payload_src2Tag;
  wire                issueQueueComponent_5_io_issueOut_payload_src2Ready;
  wire                issueQueueComponent_5_io_issueOut_payload_src2IsFpr;
  wire                issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_valid;
  wire                issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isDiv;
  wire                issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isSigned;
  wire                issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isWordOp;
  wire                issueQueueComponent_6_io_allocateIn_ready;
  wire                issueQueueComponent_6_io_issueOut_valid;
  wire       [3:0]    issueQueueComponent_6_io_issueOut_payload_robPtr;
  wire       [5:0]    issueQueueComponent_6_io_issueOut_payload_physDest_idx;
  wire                issueQueueComponent_6_io_issueOut_payload_physDestIsFpr;
  wire                issueQueueComponent_6_io_issueOut_payload_writesToPhysReg;
  wire                issueQueueComponent_6_io_issueOut_payload_useSrc1;
  wire       [31:0]   issueQueueComponent_6_io_issueOut_payload_src1Data;
  wire       [5:0]    issueQueueComponent_6_io_issueOut_payload_src1Tag;
  wire                issueQueueComponent_6_io_issueOut_payload_src1Ready;
  wire                issueQueueComponent_6_io_issueOut_payload_src1IsFpr;
  wire                issueQueueComponent_6_io_issueOut_payload_useSrc2;
  wire       [31:0]   issueQueueComponent_6_io_issueOut_payload_src2Data;
  wire       [5:0]    issueQueueComponent_6_io_issueOut_payload_src2Tag;
  wire                issueQueueComponent_6_io_issueOut_payload_src2Ready;
  wire                issueQueueComponent_6_io_issueOut_payload_src2IsFpr;
  wire       [4:0]    issueQueueComponent_6_io_issueOut_payload_branchCtrl_condition;
  wire                issueQueueComponent_6_io_issueOut_payload_branchCtrl_isJump;
  wire                issueQueueComponent_6_io_issueOut_payload_branchCtrl_isLink;
  wire       [4:0]    issueQueueComponent_6_io_issueOut_payload_branchCtrl_linkReg_idx;
  wire       [1:0]    issueQueueComponent_6_io_issueOut_payload_branchCtrl_linkReg_rtype;
  wire                issueQueueComponent_6_io_issueOut_payload_branchCtrl_isIndirect;
  wire       [2:0]    issueQueueComponent_6_io_issueOut_payload_branchCtrl_laCfIdx;
  wire       [31:0]   issueQueueComponent_6_io_issueOut_payload_imm;
  wire       [31:0]   issueQueueComponent_6_io_issueOut_payload_pc;
  wire                issueQueueComponent_6_io_issueOut_payload_branchPrediction_isTaken;
  wire       [31:0]   issueQueueComponent_6_io_issueOut_payload_branchPrediction_target;
  wire                issueQueueComponent_6_io_issueOut_payload_branchPrediction_wasPredicted;
  wire                issueQueueComponent_7_io_allocateIn_ready;
  wire                issueQueueComponent_7_io_issueOut_valid;
  wire       [3:0]    issueQueueComponent_7_io_issueOut_payload_robPtr;
  wire       [5:0]    issueQueueComponent_7_io_issueOut_payload_physDest_idx;
  wire                issueQueueComponent_7_io_issueOut_payload_physDestIsFpr;
  wire                issueQueueComponent_7_io_issueOut_payload_writesToPhysReg;
  wire                issueQueueComponent_7_io_issueOut_payload_useSrc1;
  wire       [31:0]   issueQueueComponent_7_io_issueOut_payload_src1Data;
  wire       [5:0]    issueQueueComponent_7_io_issueOut_payload_src1Tag;
  wire                issueQueueComponent_7_io_issueOut_payload_src1Ready;
  wire                issueQueueComponent_7_io_issueOut_payload_src1IsFpr;
  wire                issueQueueComponent_7_io_issueOut_payload_useSrc2;
  wire       [31:0]   issueQueueComponent_7_io_issueOut_payload_src2Data;
  wire       [5:0]    issueQueueComponent_7_io_issueOut_payload_src2Tag;
  wire                issueQueueComponent_7_io_issueOut_payload_src2Ready;
  wire                issueQueueComponent_7_io_issueOut_payload_src2IsFpr;
  wire       [1:0]    issueQueueComponent_7_io_issueOut_payload_memCtrl_size;
  wire                issueQueueComponent_7_io_issueOut_payload_memCtrl_isSignedLoad;
  wire                issueQueueComponent_7_io_issueOut_payload_memCtrl_isStore;
  wire                issueQueueComponent_7_io_issueOut_payload_memCtrl_isLoadLinked;
  wire                issueQueueComponent_7_io_issueOut_payload_memCtrl_isStoreCond;
  wire       [4:0]    issueQueueComponent_7_io_issueOut_payload_memCtrl_atomicOp;
  wire                issueQueueComponent_7_io_issueOut_payload_memCtrl_isFence;
  wire       [7:0]    issueQueueComponent_7_io_issueOut_payload_memCtrl_fenceMode;
  wire                issueQueueComponent_7_io_issueOut_payload_memCtrl_isCacheOp;
  wire       [4:0]    issueQueueComponent_7_io_issueOut_payload_memCtrl_cacheOpType;
  wire                issueQueueComponent_7_io_issueOut_payload_memCtrl_isPrefetch;
  wire       [31:0]   issueQueueComponent_7_io_issueOut_payload_imm;
  wire                issueQueueComponent_7_io_issueOut_payload_usePc;
  wire       [31:0]   issueQueueComponent_7_io_issueOut_payload_pcData;
  wire                oneShot_20_io_pulseOut;
  wire                DebugDisplayPlugin_logic_displayArea_divider_io_tick;
  wire                oneShot_21_io_pulseOut;
  wire       [63:0]   multiplierBlackbox_P;
  wire                oneShot_22_io_pulseOut;
  wire                oneShot_23_io_pulseOut;
  wire                streamDemux_1_io_input_ready;
  wire                streamDemux_1_io_outputs_0_valid;
  wire       [2:0]    streamDemux_1_io_outputs_0_payload_qPtr;
  wire       [31:0]   streamDemux_1_io_outputs_0_payload_address;
  wire                streamDemux_1_io_outputs_0_payload_alignException;
  wire       [1:0]    streamDemux_1_io_outputs_0_payload_accessSize;
  wire       [3:0]    streamDemux_1_io_outputs_0_payload_storeMask;
  wire       [5:0]    streamDemux_1_io_outputs_0_payload_basePhysReg;
  wire       [31:0]   streamDemux_1_io_outputs_0_payload_immediate;
  wire                streamDemux_1_io_outputs_0_payload_usePc;
  wire       [31:0]   streamDemux_1_io_outputs_0_payload_pc;
  wire       [3:0]    streamDemux_1_io_outputs_0_payload_robPtr;
  wire                streamDemux_1_io_outputs_0_payload_isLoad;
  wire                streamDemux_1_io_outputs_0_payload_isStore;
  wire       [5:0]    streamDemux_1_io_outputs_0_payload_physDst;
  wire       [31:0]   streamDemux_1_io_outputs_0_payload_storeData;
  wire                streamDemux_1_io_outputs_0_payload_isFlush;
  wire                streamDemux_1_io_outputs_0_payload_isIO;
  wire                streamDemux_1_io_outputs_1_valid;
  wire       [2:0]    streamDemux_1_io_outputs_1_payload_qPtr;
  wire       [31:0]   streamDemux_1_io_outputs_1_payload_address;
  wire                streamDemux_1_io_outputs_1_payload_alignException;
  wire       [1:0]    streamDemux_1_io_outputs_1_payload_accessSize;
  wire       [3:0]    streamDemux_1_io_outputs_1_payload_storeMask;
  wire       [5:0]    streamDemux_1_io_outputs_1_payload_basePhysReg;
  wire       [31:0]   streamDemux_1_io_outputs_1_payload_immediate;
  wire                streamDemux_1_io_outputs_1_payload_usePc;
  wire       [31:0]   streamDemux_1_io_outputs_1_payload_pc;
  wire       [3:0]    streamDemux_1_io_outputs_1_payload_robPtr;
  wire                streamDemux_1_io_outputs_1_payload_isLoad;
  wire                streamDemux_1_io_outputs_1_payload_isStore;
  wire       [5:0]    streamDemux_1_io_outputs_1_payload_physDst;
  wire       [31:0]   streamDemux_1_io_outputs_1_payload_storeData;
  wire                streamDemux_1_io_outputs_1_payload_isFlush;
  wire                streamDemux_1_io_outputs_1_payload_isIO;
  wire                oneShot_24_io_pulseOut;
  wire                streamArbiter_9_io_inputs_0_ready;
  wire                streamArbiter_9_io_output_valid;
  wire       [3:0]    streamArbiter_9_io_output_payload_robPtr;
  wire       [5:0]    streamArbiter_9_io_output_payload_pdest;
  wire       [31:0]   streamArbiter_9_io_output_payload_address;
  wire                streamArbiter_9_io_output_payload_isIO;
  wire       [1:0]    streamArbiter_9_io_output_payload_size;
  wire                streamArbiter_9_io_output_payload_hasEarlyException;
  wire       [7:0]    streamArbiter_9_io_output_payload_earlyExceptionCode;
  wire       [0:0]    streamArbiter_9_io_chosenOH;
  wire                oneShot_25_io_pulseOut;
  wire                FetchPipelinePlugin_logic_dispatcher_io_fetchGroupIn_ready;
  wire                FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_valid;
  wire       [31:0]   FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_pc;
  wire       [31:0]   FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_instruction;
  wire                FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isBranch;
  wire                FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isJump;
  wire                FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_jumpOffset;
  wire                FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isIdle;
  wire                FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_isTaken;
  wire       [31:0]   FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_target;
  wire                FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_wasPredicted;
  wire                FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_valid;
  wire       [31:0]   FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_payload_pc;
  wire       [2:0]    FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_payload_transactionId;
  wire                FetchPipelinePlugin_logic_dispatcher_io_softRedirect_valid;
  wire       [31:0]   FetchPipelinePlugin_logic_dispatcher_io_softRedirect_payload;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_ready;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_valid;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_pc;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_0;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_1;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_2;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_3;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isBranch;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isJump;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_jumpOffset;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isIdle;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isBranch;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isJump;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_jumpOffset;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isIdle;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isBranch;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isJump;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_jumpOffset;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isIdle;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isBranch;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isJump;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_jumpOffset;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isIdle;
  wire       [3:0]    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_branchMask;
  wire                FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_fault;
  wire       [2:0]    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_numValidInstructions;
  wire       [1:0]    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_startInstructionIndex;
  wire       [1:0]    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_occupancy;
  wire       [1:0]    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_availability;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isBranch;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isJump;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_jumpOffset;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isIdle;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isBranch;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isJump;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_jumpOffset;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isIdle;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isBranch;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isJump;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_jumpOffset;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isIdle;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isBranch;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isJump;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isDirectJump;
  wire       [31:0]   FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_jumpOffset;
  wire                FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isIdle;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_cmd_ready;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_payload_data;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_payload_error;
  wire       [3:0]    CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_payload_id;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_write_cmd_ready;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_write_rsp_valid;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_write_rsp_payload_error;
  wire       [3:0]    CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_write_rsp_payload_id;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_burst;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_burst;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_strb;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_last;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_axiOut_r_ready;
  wire                CoreMemSysPlugin_logic_readBridges_0_io_axiOut_b_ready;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_cmd_ready;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_rsp_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_rsp_payload_data;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_rsp_payload_error;
  wire       [3:0]    CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_rsp_payload_id;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_cmd_ready;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_valid;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_payload_error;
  wire       [3:0]    CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_payload_id;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_burst;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_burst;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_strb;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_last;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_r_ready;
  wire                CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_b_ready;
  wire                io_axiOut_readOnly_decoder_io_input_ar_ready;
  wire                io_axiOut_readOnly_decoder_io_input_r_valid;
  wire       [31:0]   io_axiOut_readOnly_decoder_io_input_r_payload_data;
  wire       [3:0]    io_axiOut_readOnly_decoder_io_input_r_payload_id;
  wire       [1:0]    io_axiOut_readOnly_decoder_io_input_r_payload_resp;
  wire                io_axiOut_readOnly_decoder_io_input_r_payload_last;
  wire                io_axiOut_readOnly_decoder_io_outputs_0_ar_valid;
  wire       [31:0]   io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_addr;
  wire       [3:0]    io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_id;
  wire       [7:0]    io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_len;
  wire       [2:0]    io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_size;
  wire       [1:0]    io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_burst;
  wire                io_axiOut_readOnly_decoder_io_outputs_0_r_ready;
  wire                io_axiOut_readOnly_decoder_io_outputs_1_ar_valid;
  wire       [31:0]   io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_addr;
  wire       [3:0]    io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_id;
  wire       [7:0]    io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_len;
  wire       [2:0]    io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_size;
  wire       [1:0]    io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_burst;
  wire                io_axiOut_readOnly_decoder_io_outputs_1_r_ready;
  wire                io_axiOut_readOnly_decoder_io_outputs_2_ar_valid;
  wire       [31:0]   io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_addr;
  wire       [3:0]    io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_id;
  wire       [7:0]    io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_len;
  wire       [2:0]    io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_size;
  wire       [1:0]    io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_burst;
  wire                io_axiOut_readOnly_decoder_io_outputs_2_r_ready;
  wire                io_axiOut_writeOnly_decoder_io_input_aw_ready;
  wire                io_axiOut_writeOnly_decoder_io_input_w_ready;
  wire                io_axiOut_writeOnly_decoder_io_input_b_valid;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_input_b_payload_id;
  wire       [1:0]    io_axiOut_writeOnly_decoder_io_input_b_payload_resp;
  wire                io_axiOut_writeOnly_decoder_io_outputs_0_aw_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_id;
  wire       [7:0]    io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_len;
  wire       [2:0]    io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_size;
  wire       [1:0]    io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  wire                io_axiOut_writeOnly_decoder_io_outputs_0_w_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_data;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_strb;
  wire                io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_last;
  wire                io_axiOut_writeOnly_decoder_io_outputs_0_b_ready;
  wire                io_axiOut_writeOnly_decoder_io_outputs_1_aw_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_addr;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_id;
  wire       [7:0]    io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_len;
  wire       [2:0]    io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_size;
  wire       [1:0]    io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_burst;
  wire                io_axiOut_writeOnly_decoder_io_outputs_1_w_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_data;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_strb;
  wire                io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_last;
  wire                io_axiOut_writeOnly_decoder_io_outputs_1_b_ready;
  wire                io_axiOut_writeOnly_decoder_io_outputs_2_aw_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_addr;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_id;
  wire       [7:0]    io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_len;
  wire       [2:0]    io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_size;
  wire       [1:0]    io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_burst;
  wire                io_axiOut_writeOnly_decoder_io_outputs_2_w_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_data;
  wire       [3:0]    io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_strb;
  wire                io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_last;
  wire                io_axiOut_writeOnly_decoder_io_outputs_2_b_ready;
  wire                io_axiOut_readOnly_decoder_1_io_input_ar_ready;
  wire                io_axiOut_readOnly_decoder_1_io_input_r_valid;
  wire       [31:0]   io_axiOut_readOnly_decoder_1_io_input_r_payload_data;
  wire       [3:0]    io_axiOut_readOnly_decoder_1_io_input_r_payload_id;
  wire       [1:0]    io_axiOut_readOnly_decoder_1_io_input_r_payload_resp;
  wire                io_axiOut_readOnly_decoder_1_io_input_r_payload_last;
  wire                io_axiOut_readOnly_decoder_1_io_outputs_0_ar_valid;
  wire       [31:0]   io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_addr;
  wire       [3:0]    io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_id;
  wire       [7:0]    io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_len;
  wire       [2:0]    io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_size;
  wire       [1:0]    io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_burst;
  wire                io_axiOut_readOnly_decoder_1_io_outputs_0_r_ready;
  wire                io_axiOut_readOnly_decoder_1_io_outputs_1_ar_valid;
  wire       [31:0]   io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_addr;
  wire       [3:0]    io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_id;
  wire       [7:0]    io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_len;
  wire       [2:0]    io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_size;
  wire       [1:0]    io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_burst;
  wire                io_axiOut_readOnly_decoder_1_io_outputs_1_r_ready;
  wire                io_axiOut_readOnly_decoder_1_io_outputs_2_ar_valid;
  wire       [31:0]   io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_addr;
  wire       [3:0]    io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_id;
  wire       [7:0]    io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_len;
  wire       [2:0]    io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_size;
  wire       [1:0]    io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_burst;
  wire                io_axiOut_readOnly_decoder_1_io_outputs_2_r_ready;
  wire                io_axiOut_writeOnly_decoder_1_io_input_aw_ready;
  wire                io_axiOut_writeOnly_decoder_1_io_input_w_ready;
  wire                io_axiOut_writeOnly_decoder_1_io_input_b_valid;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_input_b_payload_id;
  wire       [1:0]    io_axiOut_writeOnly_decoder_1_io_input_b_payload_resp;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_addr;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_id;
  wire       [7:0]    io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_len;
  wire       [2:0]    io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_size;
  wire       [1:0]    io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_burst;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_0_w_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_data;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_strb;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_last;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_0_b_ready;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_addr;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_id;
  wire       [7:0]    io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_len;
  wire       [2:0]    io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_size;
  wire       [1:0]    io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_burst;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_1_w_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_data;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_strb;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_last;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_1_b_ready;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_addr;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_id;
  wire       [7:0]    io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_len;
  wire       [2:0]    io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_size;
  wire       [1:0]    io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_burst;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_2_w_valid;
  wire       [31:0]   io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_data;
  wire       [3:0]    io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_strb;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_last;
  wire                io_axiOut_writeOnly_decoder_1_io_outputs_2_b_ready;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_ar_ready;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_data;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_id;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_resp;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_last;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_r_ready;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_r_ready;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_r_ready;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_aw_ready;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_w_ready;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_valid;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_payload_id;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_payload_resp;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_data;
  wire       [3:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_strb;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_last;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_b_ready;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_data;
  wire       [3:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_strb;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_last;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_b_ready;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_valid;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_data;
  wire       [3:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_strb;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_last;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_b_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_ar_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_id;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_resp;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_last;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_r_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_r_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_r_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_aw_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_w_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_valid;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_payload_id;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_payload_resp;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_strb;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_last;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_b_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_strb;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_last;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_b_ready;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_valid;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_strb;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_last;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_b_ready;
  wire                axi4ReadOnlyArbiter_3_io_inputs_0_ar_ready;
  wire                axi4ReadOnlyArbiter_3_io_inputs_0_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_resp;
  wire                axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_last;
  wire                axi4ReadOnlyArbiter_3_io_inputs_1_ar_ready;
  wire                axi4ReadOnlyArbiter_3_io_inputs_1_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_resp;
  wire                axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_last;
  wire                axi4ReadOnlyArbiter_3_io_inputs_2_ar_ready;
  wire                axi4ReadOnlyArbiter_3_io_inputs_2_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_resp;
  wire                axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_last;
  wire                axi4ReadOnlyArbiter_3_io_inputs_3_ar_ready;
  wire                axi4ReadOnlyArbiter_3_io_inputs_3_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_resp;
  wire                axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_last;
  wire                axi4ReadOnlyArbiter_3_io_output_ar_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_3_io_output_ar_payload_addr;
  wire       [6:0]    axi4ReadOnlyArbiter_3_io_output_ar_payload_id;
  wire       [7:0]    axi4ReadOnlyArbiter_3_io_output_ar_payload_len;
  wire       [2:0]    axi4ReadOnlyArbiter_3_io_output_ar_payload_size;
  wire       [1:0]    axi4ReadOnlyArbiter_3_io_output_ar_payload_burst;
  wire                axi4ReadOnlyArbiter_3_io_output_r_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_0_aw_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_0_w_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_0_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_3_io_inputs_0_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_3_io_inputs_0_b_payload_resp;
  wire                axi4WriteOnlyArbiter_3_io_inputs_1_aw_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_1_w_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_1_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_3_io_inputs_1_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_3_io_inputs_1_b_payload_resp;
  wire                axi4WriteOnlyArbiter_3_io_inputs_2_aw_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_2_w_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_2_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_3_io_inputs_2_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_3_io_inputs_2_b_payload_resp;
  wire                axi4WriteOnlyArbiter_3_io_inputs_3_aw_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_3_w_ready;
  wire                axi4WriteOnlyArbiter_3_io_inputs_3_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_3_io_inputs_3_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_3_io_inputs_3_b_payload_resp;
  wire                axi4WriteOnlyArbiter_3_io_output_aw_valid;
  wire       [31:0]   axi4WriteOnlyArbiter_3_io_output_aw_payload_addr;
  wire       [6:0]    axi4WriteOnlyArbiter_3_io_output_aw_payload_id;
  wire       [7:0]    axi4WriteOnlyArbiter_3_io_output_aw_payload_len;
  wire       [2:0]    axi4WriteOnlyArbiter_3_io_output_aw_payload_size;
  wire       [1:0]    axi4WriteOnlyArbiter_3_io_output_aw_payload_burst;
  wire                axi4WriteOnlyArbiter_3_io_output_w_valid;
  wire       [31:0]   axi4WriteOnlyArbiter_3_io_output_w_payload_data;
  wire       [3:0]    axi4WriteOnlyArbiter_3_io_output_w_payload_strb;
  wire                axi4WriteOnlyArbiter_3_io_output_w_payload_last;
  wire                axi4WriteOnlyArbiter_3_io_output_b_ready;
  wire                axi4ReadOnlyArbiter_4_io_inputs_0_ar_ready;
  wire                axi4ReadOnlyArbiter_4_io_inputs_0_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_resp;
  wire                axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_last;
  wire                axi4ReadOnlyArbiter_4_io_inputs_1_ar_ready;
  wire                axi4ReadOnlyArbiter_4_io_inputs_1_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_resp;
  wire                axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_last;
  wire                axi4ReadOnlyArbiter_4_io_inputs_2_ar_ready;
  wire                axi4ReadOnlyArbiter_4_io_inputs_2_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_resp;
  wire                axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_last;
  wire                axi4ReadOnlyArbiter_4_io_inputs_3_ar_ready;
  wire                axi4ReadOnlyArbiter_4_io_inputs_3_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_resp;
  wire                axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_last;
  wire                axi4ReadOnlyArbiter_4_io_output_ar_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_4_io_output_ar_payload_addr;
  wire       [6:0]    axi4ReadOnlyArbiter_4_io_output_ar_payload_id;
  wire       [7:0]    axi4ReadOnlyArbiter_4_io_output_ar_payload_len;
  wire       [2:0]    axi4ReadOnlyArbiter_4_io_output_ar_payload_size;
  wire       [1:0]    axi4ReadOnlyArbiter_4_io_output_ar_payload_burst;
  wire                axi4ReadOnlyArbiter_4_io_output_r_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_0_aw_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_0_w_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_0_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_4_io_inputs_0_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_4_io_inputs_0_b_payload_resp;
  wire                axi4WriteOnlyArbiter_4_io_inputs_1_aw_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_1_w_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_1_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_4_io_inputs_1_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_4_io_inputs_1_b_payload_resp;
  wire                axi4WriteOnlyArbiter_4_io_inputs_2_aw_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_2_w_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_2_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_4_io_inputs_2_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_4_io_inputs_2_b_payload_resp;
  wire                axi4WriteOnlyArbiter_4_io_inputs_3_aw_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_3_w_ready;
  wire                axi4WriteOnlyArbiter_4_io_inputs_3_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_4_io_inputs_3_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_4_io_inputs_3_b_payload_resp;
  wire                axi4WriteOnlyArbiter_4_io_output_aw_valid;
  wire       [31:0]   axi4WriteOnlyArbiter_4_io_output_aw_payload_addr;
  wire       [6:0]    axi4WriteOnlyArbiter_4_io_output_aw_payload_id;
  wire       [7:0]    axi4WriteOnlyArbiter_4_io_output_aw_payload_len;
  wire       [2:0]    axi4WriteOnlyArbiter_4_io_output_aw_payload_size;
  wire       [1:0]    axi4WriteOnlyArbiter_4_io_output_aw_payload_burst;
  wire                axi4WriteOnlyArbiter_4_io_output_w_valid;
  wire       [31:0]   axi4WriteOnlyArbiter_4_io_output_w_payload_data;
  wire       [3:0]    axi4WriteOnlyArbiter_4_io_output_w_payload_strb;
  wire                axi4WriteOnlyArbiter_4_io_output_w_payload_last;
  wire                axi4WriteOnlyArbiter_4_io_output_b_ready;
  wire                axi4ReadOnlyArbiter_5_io_inputs_0_ar_ready;
  wire                axi4ReadOnlyArbiter_5_io_inputs_0_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_resp;
  wire                axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_last;
  wire                axi4ReadOnlyArbiter_5_io_inputs_1_ar_ready;
  wire                axi4ReadOnlyArbiter_5_io_inputs_1_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_resp;
  wire                axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_last;
  wire                axi4ReadOnlyArbiter_5_io_inputs_2_ar_ready;
  wire                axi4ReadOnlyArbiter_5_io_inputs_2_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_resp;
  wire                axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_last;
  wire                axi4ReadOnlyArbiter_5_io_inputs_3_ar_ready;
  wire                axi4ReadOnlyArbiter_5_io_inputs_3_r_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_data;
  wire       [4:0]    axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_id;
  wire       [1:0]    axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_resp;
  wire                axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_last;
  wire                axi4ReadOnlyArbiter_5_io_output_ar_valid;
  wire       [31:0]   axi4ReadOnlyArbiter_5_io_output_ar_payload_addr;
  wire       [6:0]    axi4ReadOnlyArbiter_5_io_output_ar_payload_id;
  wire       [7:0]    axi4ReadOnlyArbiter_5_io_output_ar_payload_len;
  wire       [2:0]    axi4ReadOnlyArbiter_5_io_output_ar_payload_size;
  wire       [1:0]    axi4ReadOnlyArbiter_5_io_output_ar_payload_burst;
  wire                axi4ReadOnlyArbiter_5_io_output_r_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_0_aw_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_0_w_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_0_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_5_io_inputs_0_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_5_io_inputs_0_b_payload_resp;
  wire                axi4WriteOnlyArbiter_5_io_inputs_1_aw_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_1_w_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_1_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_5_io_inputs_1_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_5_io_inputs_1_b_payload_resp;
  wire                axi4WriteOnlyArbiter_5_io_inputs_2_aw_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_2_w_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_2_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_5_io_inputs_2_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_5_io_inputs_2_b_payload_resp;
  wire                axi4WriteOnlyArbiter_5_io_inputs_3_aw_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_3_w_ready;
  wire                axi4WriteOnlyArbiter_5_io_inputs_3_b_valid;
  wire       [4:0]    axi4WriteOnlyArbiter_5_io_inputs_3_b_payload_id;
  wire       [1:0]    axi4WriteOnlyArbiter_5_io_inputs_3_b_payload_resp;
  wire                axi4WriteOnlyArbiter_5_io_output_aw_valid;
  wire       [31:0]   axi4WriteOnlyArbiter_5_io_output_aw_payload_addr;
  wire       [6:0]    axi4WriteOnlyArbiter_5_io_output_aw_payload_id;
  wire       [7:0]    axi4WriteOnlyArbiter_5_io_output_aw_payload_len;
  wire       [2:0]    axi4WriteOnlyArbiter_5_io_output_aw_payload_size;
  wire       [1:0]    axi4WriteOnlyArbiter_5_io_output_aw_payload_burst;
  wire                axi4WriteOnlyArbiter_5_io_output_w_valid;
  wire       [31:0]   axi4WriteOnlyArbiter_5_io_output_w_payload_data;
  wire       [3:0]    axi4WriteOnlyArbiter_5_io_output_w_payload_strb;
  wire                axi4WriteOnlyArbiter_5_io_output_w_payload_last;
  wire                axi4WriteOnlyArbiter_5_io_output_b_ready;
  wire                io_switch_btn_buffercc_io_dataOut;
  wire       [7:0]    _zz_io_triggerIn;
  wire       [0:0]    _zz_io_triggerIn_1;
  wire       [7:0]    _zz_when_Debug_l71_13;
  wire       [7:0]    _zz_io_triggerIn_2;
  wire       [4:0]    _zz_io_triggerIn_3;
  wire       [7:0]    _zz_when_Debug_l71_1_1;
  wire       [7:0]    _zz_io_triggerIn_4;
  wire       [4:0]    _zz_io_triggerIn_5;
  wire       [7:0]    _zz_when_Debug_l71_2_1;
  wire       [7:0]    _zz_io_triggerIn_6;
  wire       [4:0]    _zz_io_triggerIn_7;
  wire       [7:0]    _zz_when_Debug_l71_3_1;
  wire       [7:0]    _zz_io_triggerIn_8;
  wire       [4:0]    _zz_io_triggerIn_9;
  wire       [7:0]    _zz_when_Debug_l71_4_1;
  reg        [0:0]    _zz_CommitPlugin_logic_s0_committedThisCycle_comb;
  wire       [0:0]    _zz_CommitPlugin_logic_s0_committedThisCycle_comb_1;
  reg        [0:0]    _zz_CommitPlugin_logic_s0_recycledThisCycle_comb;
  wire       [0:0]    _zz_CommitPlugin_logic_s0_recycledThisCycle_comb_1;
  wire       [31:0]   _zz_CommitPlugin_commitStatsReg_totalCommitted;
  wire       [31:0]   _zz_CommitPlugin_commitStatsReg_physRegRecycled;
  wire       [31:0]   _zz_CommitPlugin_commitStatsReg_robFlushCount;
  wire       [7:0]    _zz_io_triggerIn_10;
  wire       [4:0]    _zz_io_triggerIn_11;
  wire       [7:0]    _zz_when_Debug_l71_5_1;
  wire       [7:0]    _zz_io_triggerIn_12;
  wire       [4:0]    _zz_io_triggerIn_13;
  wire       [7:0]    _zz_when_Debug_l71_6_1;
  wire                _zz_DispatchPlugin_logic_dispatchOH;
  wire                _zz_DispatchPlugin_logic_dispatchOH_1;
  wire                _zz_DispatchPlugin_logic_dispatchOH_2;
  wire       [0:0]    _zz_DispatchPlugin_logic_dispatchOH_3;
  wire       [1:0]    _zz_DispatchPlugin_logic_dispatchOH_4;
  reg                 _zz_DispatchPlugin_logic_destinationIqReady_3;
  wire       [1:0]    _zz_DispatchPlugin_logic_destinationIqReady_4;
  wire       [0:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_2;
  wire       [7:0]    _zz_io_triggerIn_14;
  wire       [4:0]    _zz_io_triggerIn_15;
  wire       [7:0]    _zz_when_Debug_l71_7_1;
  wire       [63:0]   _zz_MulEU_MulEuPlugin_euResult_data_1;
  wire       [7:0]    _zz_io_triggerIn_16;
  wire       [4:0]    _zz_io_triggerIn_17;
  wire       [7:0]    _zz_when_Debug_l71_8_1;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_1;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_2;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_3;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_4;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_5;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_6;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_7;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_1;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_2;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_3;
  wire       [31:0]   _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_4;
  wire       [7:0]    _zz_io_triggerIn_18;
  wire       [4:0]    _zz_io_triggerIn_19;
  wire       [7:0]    _zz_when_Debug_l71_9_1;
  wire       [7:0]    _zz_io_triggerIn_20;
  wire       [4:0]    _zz_io_triggerIn_21;
  wire       [7:0]    _zz_when_Debug_l71_10_1;
  wire       [31:0]   _zz__zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_2;
  wire       [3:0]    _zz_LoadQueuePlugin_logic_loadQueue_pushOh;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp;
  reg        [31:0]   _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp;
  reg        [31:0]   _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp;
  wire       [2:0]    _zz_StoreBufferPlugin_logic_dcacheResponseForHead;
  wire       [7:0]    _zz_io_triggerIn_22;
  wire       [5:0]    _zz_io_triggerIn_23;
  wire       [7:0]    _zz_when_Debug_l71_11_1;
  wire       [1:0]    _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_1;
  wire       [3:0]    _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask;
  wire       [4:0]    _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_2;
  wire       [4:0]    _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_3;
  wire       [1:0]    _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_4;
  wire       [6:0]    _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_5;
  wire       [6:0]    _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_6;
  wire       [1:0]    _zz__zz_StoreBufferPlugin_logic_loadQueryBe_1;
  wire       [3:0]    _zz__zz_StoreBufferPlugin_logic_loadQueryBe;
  wire       [4:0]    _zz__zz_StoreBufferPlugin_logic_loadQueryBe_2;
  wire       [4:0]    _zz__zz_StoreBufferPlugin_logic_loadQueryBe_3;
  wire       [1:0]    _zz__zz_StoreBufferPlugin_logic_loadQueryBe_4;
  wire       [6:0]    _zz__zz_StoreBufferPlugin_logic_loadQueryBe_5;
  wire       [6:0]    _zz__zz_StoreBufferPlugin_logic_loadQueryBe_6;
  wire       [1:0]    _zz_FetchPipelinePlugin_logic_retryIdCounter_valueNext;
  wire       [0:0]    _zz_FetchPipelinePlugin_logic_retryIdCounter_valueNext_1;
  wire       [27:0]   _zz_FetchPipelinePlugin_logic_s2_logic_cmdPayload_transactionId;
  wire       [7:0]    _zz_218;
  wire       [27:0]   _zz_219;
  wire       [2:0]    _zz__zz_io_push_payload_numValidInstructions;
  reg                 _zz__zz_71;
  wire       [42:0]   _zz_ICachePlugin_logic_storage_tagLruRam_port;
  reg                 _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0;
  reg                 _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1;
  wire       [20:0]   _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag_1;
  wire       [20:0]   _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_1_tag;
  wire       [1:0]    _zz__zz_ICachePlugin_logic_pipeline_f2_hitWayIdx;
  wire       [1:0]    _zz_ICachePlugin_logic_refill_refillCounter_valueNext;
  wire       [0:0]    _zz_ICachePlugin_logic_refill_refillCounter_valueNext_1;
  wire       [127:0]  _zz_ICachePlugin_logic_storage_dataRams_0_port;
  wire       [127:0]  _zz_ICachePlugin_logic_storage_dataRams_1_port;
  wire       [9:0]    _zz_BpuPipelinePlugin_logic_pht_port;
  wire       [7:0]    _zz_BpuPipelinePlugin_logic_btb_port;
  wire       [54:0]   _zz_BpuPipelinePlugin_logic_btb_port_1;
  wire       [6:0]    _zz_io_uart_ar_bits_id;
  wire       [7:0]    _zz_uartAxi_r_payload_id;
  wire       [6:0]    _zz_io_uart_aw_bits_id;
  wire       [7:0]    _zz_uartAxi_b_payload_id;
  wire       [31:0]   _zz_io_leds_1;
  reg                 _zz_1;
  reg                 _zz_2;
  wire                BpuPipelinePlugin_logic_u2_write_ready;
  reg        [31:0]   BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_pc;
  reg                 BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken;
  reg        [31:0]   BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_target;
  wire       [31:0]   BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_pc;
  wire                BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_isTaken;
  wire       [31:0]   BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_target;
  wire                BpuPipelinePlugin_logic_u1_read_ready;
  reg        [2:0]    BpuPipelinePlugin_logic_s2_predict_TRANSACTION_ID;
  wire                BpuPipelinePlugin_logic_s2_predict_ready;
  wire       [31:0]   BpuPipelinePlugin_logic_s2_predict_TARGET_PC;
  wire                BpuPipelinePlugin_logic_s2_predict_IS_TAKEN;
  reg        [31:0]   BpuPipelinePlugin_logic_s2_predict_Q_PC;
  wire                BpuPipelinePlugin_logic_s1_read_ready;
  wire       [2:0]    BpuPipelinePlugin_logic_s1_read_TRANSACTION_ID;
  wire       [31:0]   BpuPipelinePlugin_logic_s1_read_Q_PC;
  reg                 _zz_3;
  reg                 _zz_4;
  wire                ICache_F2_HitCheck_ready;
  reg        [20:0]   ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_0_tag;
  reg        [20:0]   ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_1_tag;
  reg                 ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_lru;
  reg                 ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_USE_FORWARDED_META;
  reg                 ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_VALID_MASK_0;
  reg                 ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_VALID_MASK_1;
  reg        [31:0]   ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_address;
  reg        [7:0]    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_transactionId;
  wire       [20:0]   ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_0_tag;
  wire       [20:0]   ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_1_tag;
  wire                ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_lru;
  wire                ICache_F1_Access_ICachePlugin_logic_pipeline_F2_USE_FORWARDED_META;
  wire                ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0;
  wire                ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1;
  wire                ICache_F1_Access_ready;
  wire       [31:0]   ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_address;
  wire       [7:0]    ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_transactionId;
  wire                s4_Predecode_isFlushingRoot;
  wire                s3_ICache_Wait_isFlushingRoot;
  wire                s2_ICache_Access_isFlushingRoot;
  wire                s1_PC_Gen_isFlushingRoot;
  wire                s1_PC_Gen_isFlushed;
  wire                s2_ICache_Access_isFlushed;
  wire                s4_Predecode_isFlushed;
  wire                s3_ICache_Wait_isFlushed;
  reg        [31:0]   s2_ICache_Access_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC;
  reg        [31:0]   s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC;
  reg        [31:0]   s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC;
  reg                 s4_Predecode_ready;
  reg        [31:0]   s2_ICache_Access_FetchPipelinePlugin_logic_FetchPipeline_PC;
  wire                s2_ICache_Access_ready;
  reg                 _zz_s1_PC_Gen_haltRequest_FetchPipelinePlugin2_l381;
  reg                 s1_PC_Gen_ready;
  wire       [31:0]   s1_PC_Gen_FetchPipelinePlugin_logic_FetchPipeline_PC;
  wire       [31:0]   s1_PC_Gen_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC;
  wire                s3_Dispatch_isFlushingRoot;
  wire                s1_Rename_isFlushingRoot;
  wire                s0_Decode_isFlushingRoot;
  wire                s0_Decode_isFlushed;
  wire                s1_Rename_isFlushed;
  wire                s2_RobAlloc_isFlushed;
  wire                s3_Dispatch_isFlushed;
  wire                s3_Result_isFlushingRoot;
  wire                s2_Select_isFlushingRoot;
  wire                s1_Calc_isFlushingRoot;
  wire                s0_Dispatch_isFlushingRoot;
  wire                s0_Dispatch_isFlushed;
  wire                s1_Calc_isFlushed;
  wire                s2_Select_isFlushed;
  wire                s3_Result_isFlushed;
  wire                s3_Result_ready;
  reg        [3:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc1;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Tag;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc2;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Tag;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr;
  reg        [4:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink;
  reg        [4:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx;
  reg        [1:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect;
  reg        [2:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_imm;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_pc;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_isMispredictedBranch;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_isTaken;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_writesToPreg;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_data;
  wire                s2_Select_ready;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_data_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_data_2;
  reg        [3:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr_1;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc1_1;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data_1;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Tag_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc2_1;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data_1;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Tag_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr_1;
  reg        [4:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink_1;
  reg        [4:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx_1;
  reg        [1:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect_1;
  reg        [2:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx_1;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_1;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken_1;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted_1;
  wire                s1_Calc_ready;
  reg        [3:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr_2;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx_2;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr_2;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg_2;
  reg                 _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_valid;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data_2;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_address;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready_2;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr_2;
  reg                 _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_valid;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data_2;
  reg        [5:0]    _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_address;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready_2;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr_2;
  reg        [4:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2;
  reg                 _zz_switch_BranchEuPlugin_l133;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink_2;
  reg        [4:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx_2;
  reg        [1:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2;
  reg                 _zz_switch_BranchEuPlugin_l133_1;
  reg        [2:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx_2;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_2;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_2;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken_2;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target_2;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted_2;
  wire       [4:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3;
  wire       [1:0]    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3;
  wire       [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_3;
  wire                s0_Dispatch_ready;
  wire                mul_s7_Writeback_isFlushingRoot;
  wire                mul_s6_Execute_isFlushingRoot;
  wire                mul_s5_Execute_isFlushingRoot;
  wire                mul_s4_Execute_isFlushingRoot;
  wire                mul_s3_Execute_isFlushingRoot;
  wire                mul_s2_Execute_isFlushingRoot;
  wire                mul_s1_ReadRegs_isFlushingRoot;
  wire                mul_s0_Dispatch_isFlushingRoot;
  wire                mul_s0_Dispatch_isFlushed;
  wire                mul_s1_ReadRegs_isFlushed;
  wire                mul_s2_Execute_isFlushed;
  wire                mul_s3_Execute_isFlushed;
  wire                mul_s4_Execute_isFlushed;
  wire                mul_s5_Execute_isFlushed;
  wire                mul_s6_Execute_isFlushed;
  wire                mul_s7_Writeback_isFlushed;
  reg        [3:0]    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx;
  reg                 _zz_MulEU_MulEuPlugin_euResult_writesToPreg;
  reg                 _zz_5;
  reg                 _zz_6;
  reg                 _zz_7;
  reg        [3:0]    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_1;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_1;
  reg                 _zz_MulEU_MulEuPlugin_euResult_writesToPreg_1;
  reg                 _zz_8;
  reg                 _zz_9;
  reg                 _zz_10;
  reg        [3:0]    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_2;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_2;
  reg                 _zz_MulEU_MulEuPlugin_euResult_writesToPreg_2;
  reg                 _zz_11;
  reg                 _zz_12;
  reg                 _zz_13;
  reg        [3:0]    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_3;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_3;
  reg                 _zz_MulEU_MulEuPlugin_euResult_writesToPreg_3;
  reg                 _zz_14;
  reg                 _zz_15;
  reg                 _zz_16;
  reg        [3:0]    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_4;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_4;
  reg                 _zz_MulEU_MulEuPlugin_euResult_writesToPreg_4;
  reg                 _zz_17;
  reg                 _zz_18;
  reg                 _zz_19;
  wire                mul_s7_Writeback_ready;
  wire                mul_s2_Execute_ready;
  reg        [3:0]    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_5;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_5;
  reg                 _zz_MulEU_MulEuPlugin_euResult_writesToPreg_5;
  reg                 _zz_20;
  reg                 _zz_21;
  reg                 _zz_22;
  wire       [63:0]   _zz_MulEU_MulEuPlugin_euResult_data;
  wire       [31:0]   _zz_B;
  wire       [31:0]   _zz_A;
  wire                mul_s1_ReadRegs_ready;
  reg        [3:0]    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_6;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_6;
  reg                 _zz_MulEU_MulEuPlugin_euResult_writesToPreg_6;
  reg                 _zz_MulEU_MulEuPlugin_gprReadPorts_0_valid;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_gprReadPorts_0_address;
  reg                 _zz_MulEU_MulEuPlugin_gprReadPorts_1_valid;
  reg        [5:0]    _zz_MulEU_MulEuPlugin_gprReadPorts_1_address;
  reg                 _zz_23;
  reg                 _zz_24;
  reg                 _zz_25;
  wire                mul_s0_Dispatch_ready;
  wire                s3_Writeback_isFlushingRoot;
  wire                s2_Execute_isFlushingRoot;
  wire                s1_ReadRegs_isFlushingRoot;
  wire                s0_Dispatch_isFlushingRoot_1;
  wire                s0_Dispatch_isFlushed_1;
  wire                s1_ReadRegs_isFlushed;
  wire                s2_Execute_isFlushed;
  wire                s3_Writeback_isFlushed;
  wire                s3_Writeback_ready;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_euResult_data;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_writesToPreg;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_hasException;
  reg        [0:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode;
  reg        [3:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_robPtr;
  reg        [5:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_physDestIsFpr;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_writesToPhysReg;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_useSrc1;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data;
  reg        [5:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Tag;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Ready;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1IsFpr;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_useSrc2;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data;
  reg        [5:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Tag;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Ready;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2IsFpr;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_valid;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSub;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isAdd;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSigned;
  reg        [1:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_valid;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRight;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isArithmetic;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRotate;
  reg                 _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isDoubleWord;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_euResult_uop_imm;
  reg        [2:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage;
  wire                s2_Execute_ready;
  wire       [0:0]    _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_1;
  reg        [31:0]   _zz_io_iqEntryIn_payload_src2Data;
  reg        [31:0]   _zz_io_iqEntryIn_payload_src1Data;
  reg        [3:0]    _zz_io_iqEntryIn_payload_robPtr;
  reg        [5:0]    _zz_io_iqEntryIn_payload_physDest_idx;
  reg                 _zz_io_iqEntryIn_payload_physDestIsFpr;
  reg                 _zz_io_iqEntryIn_payload_writesToPhysReg;
  reg                 _zz_io_iqEntryIn_payload_useSrc1;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data_1;
  reg        [5:0]    _zz_io_iqEntryIn_payload_src1Tag;
  reg                 _zz_io_iqEntryIn_payload_src1Ready;
  reg                 _zz_io_iqEntryIn_payload_src1IsFpr;
  reg                 _zz_io_iqEntryIn_payload_useSrc2;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data_1;
  reg        [5:0]    _zz_io_iqEntryIn_payload_src2Tag;
  reg                 _zz_io_iqEntryIn_payload_src2Ready;
  reg                 _zz_io_iqEntryIn_payload_src2IsFpr;
  reg                 _zz_io_iqEntryIn_payload_aluCtrl_valid;
  reg                 _zz_io_iqEntryIn_payload_aluCtrl_isSub;
  reg                 _zz_io_iqEntryIn_payload_aluCtrl_isAdd;
  reg                 _zz_io_iqEntryIn_payload_aluCtrl_isSigned;
  reg        [1:0]    _zz_io_iqEntryIn_payload_aluCtrl_logicOp;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_valid;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_isRight;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_isArithmetic;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_isRotate;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_isDoubleWord;
  reg        [31:0]   _zz_io_iqEntryIn_payload_imm;
  reg        [2:0]    _zz_io_iqEntryIn_payload_immUsage;
  wire                s1_ReadRegs_ready;
  reg        [3:0]    _zz_io_iqEntryIn_payload_robPtr_1;
  reg        [5:0]    _zz_io_iqEntryIn_payload_physDest_idx_1;
  reg                 _zz_io_iqEntryIn_payload_physDestIsFpr_1;
  reg                 _zz_io_iqEntryIn_payload_writesToPhysReg_1;
  reg                 _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_valid;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data_2;
  reg        [5:0]    _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_address;
  reg                 _zz_io_iqEntryIn_payload_src1Ready_1;
  reg                 _zz_io_iqEntryIn_payload_src1IsFpr_1;
  reg                 _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_valid;
  reg        [31:0]   _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data_2;
  reg        [5:0]    _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_address;
  reg                 _zz_io_iqEntryIn_payload_src2Ready_1;
  reg                 _zz_io_iqEntryIn_payload_src2IsFpr_1;
  reg                 _zz_io_iqEntryIn_payload_aluCtrl_valid_1;
  reg                 _zz_io_iqEntryIn_payload_aluCtrl_isSub_1;
  reg                 _zz_io_iqEntryIn_payload_aluCtrl_isAdd_1;
  reg                 _zz_io_iqEntryIn_payload_aluCtrl_isSigned_1;
  reg        [1:0]    _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_valid_1;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_isRight_1;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_isArithmetic_1;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_isRotate_1;
  reg                 _zz_io_iqEntryIn_payload_shiftCtrl_isDoubleWord_1;
  reg        [31:0]   _zz_io_iqEntryIn_payload_imm_1;
  reg        [2:0]    _zz_io_iqEntryIn_payload_immUsage_1;
  wire       [1:0]    _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2;
  wire       [2:0]    _zz_io_iqEntryIn_payload_immUsage_2;
  wire                s0_Dispatch_ready_1;
  reg                 when_Connection_l66;
  wire       [31:0]   s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode;
  wire       [3:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr;
  wire       [31:0]   s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm;
  wire       [2:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence;
  wire       [7:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect;
  wire       [2:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx;
  wire       [3:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
  wire       [2:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond;
  wire       [13:0]   s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
  wire       [19:0]   s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp;
  wire       [3:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode;
  wire       [7:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken;
  wire       [31:0]   s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted;
  wire       [5:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr;
  wire       [5:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr;
  wire       [5:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr;
  wire       [5:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg;
  wire       [3:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr;
  wire       [15:0]   s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_executed;
  wire                s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException;
  wire       [7:0]    s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode;
  reg                 _zz_s1_Rename_isFlushingRoot;
  wire       [31:0]   s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_pc;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isValid;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode;
  wire       [3:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_idx;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_writeArchDestEn;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_idx;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_useArchSrc1;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_idx;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_useArchSrc2;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_usePcForAddr;
  wire       [31:0]   s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_imm;
  wire       [2:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_valid;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isSub;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isAdd;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isSigned;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_valid;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isRight;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isArithmetic;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isRotate;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_valid;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isDiv;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isSigned;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isWordOp;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isSignedLoad;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isStore;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isLoadLinked;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isStoreCond;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_atomicOp;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isFence;
  wire       [7:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_fenceMode;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isCacheOp;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_cacheOpType;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isPrefetch;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isJump;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isLink;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isIndirect;
  wire       [2:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_laCfIdx;
  wire       [3:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_opType;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
  wire       [2:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_roundingMode;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fcmpCond;
  wire       [13:0]   s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_csrAddr;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isWrite;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isRead;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isExchange;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
  wire       [19:0]   s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_sysCode;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_isTlbOp;
  wire       [3:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_tlbOpType;
  wire       [1:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_hasDecodeException;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isMicrocode;
  wire       [7:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_microcodeEntry;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isSerializing;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isBranchOrJump;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_isTaken;
  wire       [31:0]   s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_target;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_wasPredicted;
  wire       [5:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc1_idx;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc1IsFpr;
  wire       [5:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc2_idx;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc2IsFpr;
  wire       [5:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physDest_idx;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physDestIsFpr;
  wire       [5:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_oldPhysDest_idx;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_oldPhysDestIsFpr;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_allocatesPhysDest;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_writesToPhysReg;
  wire       [3:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_robPtr;
  wire       [15:0]   s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_uniqueId;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_dispatched;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_executed;
  wire                s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_hasException;
  wire       [7:0]    s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_exceptionCode;
  reg                 _zz_s2_RobAlloc_haltRequest_RenamePlugin_l85;
  reg                 s2_RobAlloc_IssuePipelineSignals_NEEDS_PHYS_REG_0;
  reg        [31:0]   s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_pc;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isValid;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode;
  reg        [3:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr;
  reg        [31:0]   s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_imm;
  reg        [2:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence;
  reg        [7:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect;
  reg        [2:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx;
  reg        [3:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest;
  reg        [2:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond;
  reg        [13:0]   s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc;
  reg        [19:0]   s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp;
  reg        [3:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType;
  reg        [1:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode;
  reg        [7:0]    s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isSerializing;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken;
  reg        [31:0]   s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target;
  reg                 s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted;
  wire                s1_Rename_IssuePipelineSignals_NEEDS_PHYS_REG_0;
  reg        [31:0]   s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_pc;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isValid;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode;
  reg        [3:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr;
  reg        [31:0]   s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_imm;
  reg        [2:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence;
  reg        [7:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect;
  reg        [2:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx;
  reg        [3:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest;
  reg        [2:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond;
  reg        [13:0]   s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc;
  reg        [19:0]   s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp;
  reg        [3:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType;
  reg        [1:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode;
  reg        [7:0]    s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isSerializing;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken;
  reg        [31:0]   s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target;
  reg                 s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted;
  reg                 _zz_s0_Decode_isFlushingRoot;
  reg        [31:0]   s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode;
  reg        [3:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr;
  reg        [31:0]   s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm;
  reg        [2:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence;
  reg        [7:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect;
  reg        [2:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode;
  reg        [7:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken;
  reg        [31:0]   s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr;
  reg        [5:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr;
  reg        [5:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr;
  reg        [5:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg;
  reg        [3:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr;
  reg        [15:0]   s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_executed;
  reg                 s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException;
  reg        [7:0]    s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode;
  reg                 s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_isTaken;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_target;
  reg                 s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_wasPredicted;
  reg                 s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_isTaken;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_target;
  reg                 s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_wasPredicted;
  reg                 s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_isTaken;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_target;
  reg                 s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_wasPredicted;
  reg                 s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_isTaken;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_target;
  reg                 s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_wasPredicted;
  wire       [31:0]   s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_pc;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isValid;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode;
  wire       [3:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr;
  wire       [31:0]   s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_imm;
  wire       [2:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence;
  wire       [7:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect;
  wire       [2:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx;
  wire       [3:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest;
  wire       [2:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond;
  wire       [13:0]   s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc;
  wire       [19:0]   s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp;
  wire       [3:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType;
  wire       [1:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode;
  wire       [7:0]    s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isSerializing;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken;
  wire       [31:0]   s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target;
  wire                s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted;
  reg        [3:0]    s0_Decode_IssuePipelineSignals_VALID_MASK;
  reg                 s0_Decode_IssuePipelineSignals_IS_FAULT_IN;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_0;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_1;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_2;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_3;
  reg        [31:0]   s0_Decode_IssuePipelineSignals_GROUP_PC_IN;
  reg                 s3_Dispatch_ready;
  reg                 s2_RobAlloc_ready;
  wire                s1_Rename_ready;
  wire                s0_Decode_ready;
  wire                BpuPipelinePlugin_queryPortIn_valid;
  wire       [31:0]   BpuPipelinePlugin_queryPortIn_payload_pc;
  wire       [2:0]    BpuPipelinePlugin_queryPortIn_payload_transactionId;
  wire                BpuPipelinePlugin_responseFlowOut_valid;
  wire                BpuPipelinePlugin_responseFlowOut_payload_isTaken;
  wire       [31:0]   BpuPipelinePlugin_responseFlowOut_payload_target;
  wire       [2:0]    BpuPipelinePlugin_responseFlowOut_payload_transactionId;
  wire       [31:0]   BpuPipelinePlugin_responseFlowOut_payload_qPc;
  reg                 BpuPipelinePlugin_updatePortIn_valid;
  wire                BpuPipelinePlugin_updatePortIn_ready;
  reg        [31:0]   BpuPipelinePlugin_updatePortIn_payload_pc;
  reg                 BpuPipelinePlugin_updatePortIn_payload_isTaken;
  reg        [31:0]   BpuPipelinePlugin_updatePortIn_payload_target;
  reg        [15:0]   FetchPipelinePlugin_dbg_cycles;
  reg        [2:0]    FetchPipelinePlugin_dbg_c;
  wire                FetchPipelinePlugin_doHardRedirect_listening;
  wire                FetchPipelinePlugin_doSoftRedirect_listening;
  wire       [63:0]   BusyTablePlugin_combinationalBusyBits;
  wire                ROBPlugin_aggregatedFlushSignal_valid;
  wire       [1:0]    ROBPlugin_aggregatedFlushSignal_payload_reason;
  wire       [3:0]    ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr;
  reg                 CheckpointManagerPlugin_saveCheckpointTrigger;
  reg                 CheckpointManagerPlugin_restoreCheckpointTrigger;
  wire                CommitPlugin_commitEnableExt;
  reg        [0:0]    CommitPlugin_commitStatsReg_committedThisCycle;
  reg        [31:0]   CommitPlugin_commitStatsReg_totalCommitted;
  reg        [31:0]   CommitPlugin_commitStatsReg_robFlushCount;
  reg        [31:0]   CommitPlugin_commitStatsReg_physRegRecycled;
  reg                 CommitPlugin_commitStatsReg_commitOOB;
  reg        [31:0]   CommitPlugin_commitStatsReg_maxCommitPc;
  wire       [31:0]   CommitPlugin_maxCommitPcExt;
  wire                CommitPlugin_maxCommitPcEnabledExt;
  (* mark_debug = "true" *) reg        [31:0]   CommitPlugin_maxCommitPcReg;
  (* mark_debug = "true" *) reg                 CommitPlugin_commitOOBReg;
  reg                 AluIntEU_AluIntEuPlugin_euResult_valid;
  reg        [3:0]    AluIntEU_AluIntEuPlugin_euResult_uop_robPtr;
  reg        [5:0]    AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_physDestIsFpr;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_writesToPhysReg;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_useSrc1;
  reg        [31:0]   AluIntEU_AluIntEuPlugin_euResult_uop_src1Data;
  reg        [5:0]    AluIntEU_AluIntEuPlugin_euResult_uop_src1Tag;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_src1Ready;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_src1IsFpr;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_useSrc2;
  reg        [31:0]   AluIntEU_AluIntEuPlugin_euResult_uop_src2Data;
  reg        [5:0]    AluIntEU_AluIntEuPlugin_euResult_uop_src2Tag;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_src2Ready;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_src2IsFpr;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_valid;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSub;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isAdd;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSigned;
  reg        [1:0]    AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_valid;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRight;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isArithmetic;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRotate;
  reg                 AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isDoubleWord;
  reg        [31:0]   AluIntEU_AluIntEuPlugin_euResult_uop_imm;
  reg        [2:0]    AluIntEU_AluIntEuPlugin_euResult_uop_immUsage;
  reg        [31:0]   AluIntEU_AluIntEuPlugin_euResult_data;
  reg                 AluIntEU_AluIntEuPlugin_euResult_writesToPreg;
  wire                AluIntEU_AluIntEuPlugin_euResult_isMispredictedBranch;
  wire                AluIntEU_AluIntEuPlugin_euResult_isTaken;
  reg                 AluIntEU_AluIntEuPlugin_euResult_hasException;
  reg        [7:0]    AluIntEU_AluIntEuPlugin_euResult_exceptionCode;
  reg                 AluIntEU_AluIntEuPlugin_euResult_destIsFpr;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_0_0_0;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_0_0_1;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_0_0_2;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_0_0_3;
  reg                 MulEU_MulEuPlugin_euResult_valid;
  wire       [31:0]   MulEU_MulEuPlugin_euResult_uop_uop_decoded_pc;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_isValid;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode;
  wire       [3:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_idx;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_writeArchDestEn;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_idx;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_useArchSrc1;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_idx;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_useArchSrc2;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_usePcForAddr;
  wire       [31:0]   MulEU_MulEuPlugin_euResult_uop_uop_decoded_imm;
  wire       [2:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_valid;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_isSub;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_isAdd;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_isSigned;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_valid;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_isRight;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_isArithmetic;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_isRotate;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_isDoubleWord;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_mulDivCtrl_valid;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_mulDivCtrl_isDiv;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_mulDivCtrl_isSigned;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_mulDivCtrl_isWordOp;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isSignedLoad;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isStore;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isLoadLinked;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isStoreCond;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_atomicOp;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isFence;
  wire       [7:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_fenceMode;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isCacheOp;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_cacheOpType;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isPrefetch;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_isJump;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_isLink;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_isIndirect;
  wire       [2:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_laCfIdx;
  wire       [3:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_opType;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest;
  wire       [2:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_roundingMode;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_isIntegerDest;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_isSignedCvt;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fcmpCond;
  wire       [13:0]   MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_csrAddr;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_isWrite;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_isRead;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_isExchange;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_useUimmAsSrc;
  wire       [19:0]   MulEU_MulEuPlugin_euResult_uop_uop_decoded_sysCtrl_sysCode;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_sysCtrl_isExceptionReturn;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_sysCtrl_isTlbOp;
  wire       [3:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_sysCtrl_tlbOpType;
  wire       [1:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_hasDecodeException;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_isMicrocode;
  wire       [7:0]    MulEU_MulEuPlugin_euResult_uop_uop_decoded_microcodeEntry;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_isSerializing;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_isBranchOrJump;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchPrediction_isTaken;
  wire       [31:0]   MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchPrediction_target;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchPrediction_wasPredicted;
  wire       [5:0]    MulEU_MulEuPlugin_euResult_uop_uop_rename_physSrc1_idx;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_rename_physSrc1IsFpr;
  wire       [5:0]    MulEU_MulEuPlugin_euResult_uop_uop_rename_physSrc2_idx;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_rename_physSrc2IsFpr;
  wire       [5:0]    MulEU_MulEuPlugin_euResult_uop_uop_rename_physDest_idx;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_rename_physDestIsFpr;
  wire       [5:0]    MulEU_MulEuPlugin_euResult_uop_uop_rename_oldPhysDest_idx;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_rename_oldPhysDestIsFpr;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_rename_allocatesPhysDest;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_rename_writesToPhysReg;
  wire       [3:0]    MulEU_MulEuPlugin_euResult_uop_uop_robPtr;
  wire       [15:0]   MulEU_MulEuPlugin_euResult_uop_uop_uniqueId;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_dispatched;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_executed;
  wire                MulEU_MulEuPlugin_euResult_uop_uop_hasException;
  wire       [7:0]    MulEU_MulEuPlugin_euResult_uop_uop_exceptionCode;
  reg        [3:0]    MulEU_MulEuPlugin_euResult_uop_robPtr;
  reg        [5:0]    MulEU_MulEuPlugin_euResult_uop_physDest_idx;
  wire                MulEU_MulEuPlugin_euResult_uop_physDestIsFpr;
  wire                MulEU_MulEuPlugin_euResult_uop_writesToPhysReg;
  wire                MulEU_MulEuPlugin_euResult_uop_useSrc1;
  wire       [31:0]   MulEU_MulEuPlugin_euResult_uop_src1Data;
  wire       [5:0]    MulEU_MulEuPlugin_euResult_uop_src1Tag;
  wire                MulEU_MulEuPlugin_euResult_uop_src1Ready;
  wire                MulEU_MulEuPlugin_euResult_uop_src1IsFpr;
  wire                MulEU_MulEuPlugin_euResult_uop_useSrc2;
  wire       [31:0]   MulEU_MulEuPlugin_euResult_uop_src2Data;
  wire       [5:0]    MulEU_MulEuPlugin_euResult_uop_src2Tag;
  wire                MulEU_MulEuPlugin_euResult_uop_src2Ready;
  wire                MulEU_MulEuPlugin_euResult_uop_src2IsFpr;
  wire                MulEU_MulEuPlugin_euResult_uop_mulDivCtrl_valid;
  wire                MulEU_MulEuPlugin_euResult_uop_mulDivCtrl_isDiv;
  wire                MulEU_MulEuPlugin_euResult_uop_mulDivCtrl_isSigned;
  wire                MulEU_MulEuPlugin_euResult_uop_mulDivCtrl_isWordOp;
  reg        [31:0]   MulEU_MulEuPlugin_euResult_data;
  reg                 MulEU_MulEuPlugin_euResult_writesToPreg;
  wire                MulEU_MulEuPlugin_euResult_isMispredictedBranch;
  wire                MulEU_MulEuPlugin_euResult_isTaken;
  reg                 MulEU_MulEuPlugin_euResult_hasException;
  reg        [7:0]    MulEU_MulEuPlugin_euResult_exceptionCode;
  reg                 MulEU_MulEuPlugin_euResult_destIsFpr;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_1_0_0;
  reg                 BranchEU_BranchEuPlugin_euResult_valid;
  reg        [3:0]    BranchEU_BranchEuPlugin_euResult_uop_robPtr;
  reg        [5:0]    BranchEU_BranchEuPlugin_euResult_uop_physDest_idx;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_useSrc1;
  reg        [31:0]   BranchEU_BranchEuPlugin_euResult_uop_src1Data;
  reg        [5:0]    BranchEU_BranchEuPlugin_euResult_uop_src1Tag;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_src1Ready;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_useSrc2;
  reg        [31:0]   BranchEU_BranchEuPlugin_euResult_uop_src2Data;
  reg        [5:0]    BranchEU_BranchEuPlugin_euResult_uop_src2Tag;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_src2Ready;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr;
  reg        [4:0]    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink;
  reg        [4:0]    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx;
  reg        [1:0]    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect;
  reg        [2:0]    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx;
  reg        [31:0]   BranchEU_BranchEuPlugin_euResult_uop_imm;
  reg        [31:0]   BranchEU_BranchEuPlugin_euResult_uop_pc;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken;
  reg        [31:0]   BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target;
  reg                 BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted;
  reg        [31:0]   BranchEU_BranchEuPlugin_euResult_data;
  reg                 BranchEU_BranchEuPlugin_euResult_writesToPreg;
  reg                 BranchEU_BranchEuPlugin_euResult_isMispredictedBranch;
  reg                 BranchEU_BranchEuPlugin_euResult_isTaken;
  reg                 BranchEU_BranchEuPlugin_euResult_hasException;
  reg        [7:0]    BranchEU_BranchEuPlugin_euResult_exceptionCode;
  reg                 BranchEU_BranchEuPlugin_euResult_destIsFpr;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_2_0_0;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_2_0_1;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_2_0_2;
  reg                 LsuEU_LsuEuPlugin_euResult_valid;
  reg        [3:0]    LsuEU_LsuEuPlugin_euResult_uop_robPtr;
  reg        [5:0]    LsuEU_LsuEuPlugin_euResult_uop_physDest_idx;
  wire                LsuEU_LsuEuPlugin_euResult_uop_physDestIsFpr;
  reg                 LsuEU_LsuEuPlugin_euResult_uop_writesToPhysReg;
  wire                LsuEU_LsuEuPlugin_euResult_uop_useSrc1;
  wire       [31:0]   LsuEU_LsuEuPlugin_euResult_uop_src1Data;
  wire       [5:0]    LsuEU_LsuEuPlugin_euResult_uop_src1Tag;
  wire                LsuEU_LsuEuPlugin_euResult_uop_src1Ready;
  wire                LsuEU_LsuEuPlugin_euResult_uop_src1IsFpr;
  wire                LsuEU_LsuEuPlugin_euResult_uop_useSrc2;
  wire       [31:0]   LsuEU_LsuEuPlugin_euResult_uop_src2Data;
  wire       [5:0]    LsuEU_LsuEuPlugin_euResult_uop_src2Tag;
  wire                LsuEU_LsuEuPlugin_euResult_uop_src2Ready;
  wire                LsuEU_LsuEuPlugin_euResult_uop_src2IsFpr;
  wire       [1:0]    LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size;
  wire                LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isSignedLoad;
  wire                LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isStore;
  wire                LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isLoadLinked;
  wire                LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isStoreCond;
  wire       [4:0]    LsuEU_LsuEuPlugin_euResult_uop_memCtrl_atomicOp;
  wire                LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isFence;
  wire       [7:0]    LsuEU_LsuEuPlugin_euResult_uop_memCtrl_fenceMode;
  wire                LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isCacheOp;
  wire       [4:0]    LsuEU_LsuEuPlugin_euResult_uop_memCtrl_cacheOpType;
  wire                LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isPrefetch;
  wire       [31:0]   LsuEU_LsuEuPlugin_euResult_uop_imm;
  wire                LsuEU_LsuEuPlugin_euResult_uop_usePc;
  wire       [31:0]   LsuEU_LsuEuPlugin_euResult_uop_pcData;
  wire       [31:0]   LsuEU_LsuEuPlugin_euResult_data;
  reg                 LsuEU_LsuEuPlugin_euResult_writesToPreg;
  wire                LsuEU_LsuEuPlugin_euResult_isMispredictedBranch;
  wire                LsuEU_LsuEuPlugin_euResult_isTaken;
  reg                 LsuEU_LsuEuPlugin_euResult_hasException;
  reg        [7:0]    LsuEU_LsuEuPlugin_euResult_exceptionCode;
  reg                 LsuEU_LsuEuPlugin_euResult_destIsFpr;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_3_0_0;
  wire       [4:0]    DispatchPlugin_logic_iqRegs_3_0_1;
  wire                ICachePlugin_port_cmd_valid;
  wire       [31:0]   ICachePlugin_port_cmd_payload_address;
  wire       [7:0]    ICachePlugin_port_cmd_payload_transactionId;
  reg                 ICachePlugin_port_rsp_valid;
  reg        [7:0]    ICachePlugin_port_rsp_payload_transactionId;
  reg        [31:0]   ICachePlugin_port_rsp_payload_instructions_0;
  reg        [31:0]   ICachePlugin_port_rsp_payload_instructions_1;
  reg        [31:0]   ICachePlugin_port_rsp_payload_instructions_2;
  reg        [31:0]   ICachePlugin_port_rsp_payload_instructions_3;
  reg                 ICachePlugin_port_rsp_payload_wasHit;
  reg                 ICachePlugin_port_rsp_payload_redo;
  wire                ICachePlugin_invalidate;
  reg        [7:0]    _zz_when_Debug_l71;
  wire                DataCachePlugin_setup_writebackBusy;
  wire       [7:0]    DataCachePlugin_setup_refillCompletions;
  wire                DataCachePlugin_setup_dcacheMaster_aw_valid;
  wire                DataCachePlugin_setup_dcacheMaster_aw_ready;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_aw_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_aw_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_aw_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_aw_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_aw_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_aw_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_w_valid;
  wire                DataCachePlugin_setup_dcacheMaster_w_ready;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_w_payload_data;
  wire       [3:0]    DataCachePlugin_setup_dcacheMaster_w_payload_strb;
  wire                DataCachePlugin_setup_dcacheMaster_w_payload_last;
  wire                DataCachePlugin_setup_dcacheMaster_b_valid;
  reg                 DataCachePlugin_setup_dcacheMaster_b_ready;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_b_payload_id;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_b_payload_resp;
  wire                DataCachePlugin_setup_dcacheMaster_ar_valid;
  wire                DataCachePlugin_setup_dcacheMaster_ar_ready;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_ar_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_ar_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_ar_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_ar_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_ar_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_ar_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_r_valid;
  reg                 DataCachePlugin_setup_dcacheMaster_r_ready;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_r_payload_data;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_r_payload_id;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_r_payload_resp;
  wire                DataCachePlugin_setup_dcacheMaster_r_payload_last;
  wire                io_mem_toAxi4_arCmdStaged_valid;
  wire                io_mem_toAxi4_arCmdStaged_ready;
  wire       [2:0]    io_mem_toAxi4_arCmdStaged_payload_id;
  wire       [31:0]   io_mem_toAxi4_arCmdStaged_payload_address;
  reg                 io_mem_read_cmd_rValid;
  reg        [2:0]    io_mem_read_cmd_rData_id;
  reg        [31:0]   io_mem_read_cmd_rData_address;
  wire                when_Stream_l477;
  wire                io_mem_toAxi4_rRspStaged_valid;
  wire                io_mem_toAxi4_rRspStaged_ready;
  wire       [31:0]   io_mem_toAxi4_rRspStaged_payload_data;
  wire       [2:0]    io_mem_toAxi4_rRspStaged_payload_id;
  wire       [1:0]    io_mem_toAxi4_rRspStaged_payload_resp;
  wire                io_mem_toAxi4_rRspStaged_payload_last;
  reg                 DataCachePlugin_setup_dcacheMaster_r_rValid;
  reg        [31:0]   DataCachePlugin_setup_dcacheMaster_r_rData_data;
  reg        [2:0]    DataCachePlugin_setup_dcacheMaster_r_rData_id;
  reg        [1:0]    DataCachePlugin_setup_dcacheMaster_r_rData_resp;
  reg                 DataCachePlugin_setup_dcacheMaster_r_rData_last;
  wire                when_Stream_l477_1;
  wire                io_mem_toAxi4_awRaw_valid;
  reg                 io_mem_toAxi4_awRaw_ready;
  wire                io_mem_toAxi4_awRaw_payload_last;
  wire       [31:0]   io_mem_toAxi4_awRaw_payload_fragment_address;
  wire       [31:0]   io_mem_toAxi4_awRaw_payload_fragment_data;
  wire       [2:0]    io_mem_toAxi4_awRaw_payload_fragment_id;
  wire                io_mem_toAxi4_wRaw_valid;
  wire                io_mem_toAxi4_wRaw_ready;
  wire                io_mem_toAxi4_wRaw_payload_last;
  wire       [31:0]   io_mem_toAxi4_wRaw_payload_fragment_address;
  wire       [31:0]   io_mem_toAxi4_wRaw_payload_fragment_data;
  wire       [2:0]    io_mem_toAxi4_wRaw_payload_fragment_id;
  reg                 io_mem_write_cmd_fork2_logic_linkEnable_0;
  reg                 io_mem_write_cmd_fork2_logic_linkEnable_1;
  wire                when_Stream_l1253;
  wire                when_Stream_l1253_1;
  wire                io_mem_toAxi4_awRaw_fire;
  wire                io_mem_toAxi4_wRaw_fire;
  reg                 io_mem_toAxi4_awRaw_payload_first;
  wire                when_Stream_l581;
  reg                 io_mem_toAxi4_awFiltred_valid;
  reg                 io_mem_toAxi4_awFiltred_ready;
  wire                io_mem_toAxi4_awFiltred_payload_last;
  wire       [31:0]   io_mem_toAxi4_awFiltred_payload_fragment_address;
  wire       [31:0]   io_mem_toAxi4_awFiltred_payload_fragment_data;
  wire       [2:0]    io_mem_toAxi4_awFiltred_payload_fragment_id;
  wire                io_mem_toAxi4_aw_valid;
  wire                io_mem_toAxi4_aw_ready;
  wire                io_mem_toAxi4_aw_payload_last;
  wire       [31:0]   io_mem_toAxi4_aw_payload_fragment_address;
  wire       [31:0]   io_mem_toAxi4_aw_payload_fragment_data;
  wire       [2:0]    io_mem_toAxi4_aw_payload_fragment_id;
  reg                 io_mem_toAxi4_awFiltred_rValid;
  reg                 io_mem_toAxi4_awFiltred_rData_last;
  reg        [31:0]   io_mem_toAxi4_awFiltred_rData_fragment_address;
  reg        [31:0]   io_mem_toAxi4_awFiltred_rData_fragment_data;
  reg        [2:0]    io_mem_toAxi4_awFiltred_rData_fragment_id;
  wire                when_Stream_l477_2;
  wire                _zz_io_mem_toAxi4_wRaw_ready;
  wire                io_mem_toAxi4_w_valid;
  reg                 io_mem_toAxi4_w_ready;
  wire                io_mem_toAxi4_w_payload_last;
  wire       [31:0]   io_mem_toAxi4_w_payload_fragment_address;
  wire       [31:0]   io_mem_toAxi4_w_payload_fragment_data;
  wire       [2:0]    io_mem_toAxi4_w_payload_fragment_id;
  wire                io_mem_toAxi4_wStaged_valid;
  wire                io_mem_toAxi4_wStaged_ready;
  wire                io_mem_toAxi4_wStaged_payload_last;
  wire       [31:0]   io_mem_toAxi4_wStaged_payload_fragment_address;
  wire       [31:0]   io_mem_toAxi4_wStaged_payload_fragment_data;
  wire       [2:0]    io_mem_toAxi4_wStaged_payload_fragment_id;
  reg                 io_mem_toAxi4_w_rValid;
  reg                 io_mem_toAxi4_w_rData_last;
  reg        [31:0]   io_mem_toAxi4_w_rData_fragment_address;
  reg        [31:0]   io_mem_toAxi4_w_rData_fragment_data;
  reg        [2:0]    io_mem_toAxi4_w_rData_fragment_id;
  wire                when_Stream_l477_3;
  wire                io_mem_toAxi4_bRspStaged_valid;
  wire                io_mem_toAxi4_bRspStaged_ready;
  wire       [2:0]    io_mem_toAxi4_bRspStaged_payload_id;
  wire       [1:0]    io_mem_toAxi4_bRspStaged_payload_resp;
  reg                 DataCachePlugin_setup_dcacheMaster_b_rValid;
  reg        [2:0]    DataCachePlugin_setup_dcacheMaster_b_rData_id;
  reg        [1:0]    DataCachePlugin_setup_dcacheMaster_b_rData_resp;
  wire                when_Stream_l477_4;
  wire       [0:0]    _zz_when_Debug_l71_1;
  wire                when_Debug_l71;
  reg        [63:0]   BusyTablePlugin_early_setup_busyTableReg;
  reg        [63:0]   BusyTablePlugin_early_setup_clearMask;
  reg        [63:0]   BusyTablePlugin_early_setup_setMask;
  wire                s0_Decode_valid;
  reg                 _zz_s1_Rename_valid;
  reg                 s1_Rename_valid;
  reg                 _zz_s2_RobAlloc_valid;
  reg                 s2_RobAlloc_valid;
  reg                 _zz_s3_Dispatch_valid;
  reg                 s3_Dispatch_valid;
  wire                s0_Decode_isFiring;
  wire       [4:0]    _zz_when_Debug_l71_2;
  wire                when_Debug_l71_1;
  wire                s1_Rename_isFiring;
  wire       [4:0]    _zz_when_Debug_l71_3;
  wire                when_Debug_l71_2;
  wire                s2_RobAlloc_isFiring;
  wire       [4:0]    _zz_when_Debug_l71_4;
  wire                when_Debug_l71_3;
  wire                s3_Dispatch_isFiring;
  wire       [4:0]    _zz_when_Debug_l71_5;
  wire                when_Debug_l71_4;
  reg                 CommitPlugin_hw_busyTableClearPort_valid;
  reg        [5:0]    CommitPlugin_hw_busyTableClearPort_payload;
  reg                 CommitPlugin_hw_robFlushPort_valid;
  reg        [1:0]    CommitPlugin_hw_robFlushPort_payload_reason;
  reg        [3:0]    CommitPlugin_hw_robFlushPort_payload_targetRobPtr;
  reg                 CommitPlugin_hw_redirectPort_valid;
  reg        [31:0]   CommitPlugin_hw_redirectPort_payload;
  wire                RenamePlugin_setup_btSetBusyPorts_0_valid;
  wire       [5:0]    RenamePlugin_setup_btSetBusyPorts_0_payload;
  wire                AluIntEU_AluIntEuPlugin_wakeupSourcePort_valid;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_wakeupSourcePort_payload_physRegIdx;
  wire                AluIntEU_AluIntEuPlugin_gprReadPorts_0_valid;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_gprReadPorts_0_address;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp;
  wire                AluIntEU_AluIntEuPlugin_gprReadPorts_1_valid;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_gprReadPorts_1_address;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp;
  wire                AluIntEU_AluIntEuPlugin_gprWritePort_valid;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_gprWritePort_address;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_gprWritePort_data;
  wire                AluIntEU_AluIntEuPlugin_bypassOutputPort_valid;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_physRegIdx;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_physRegData;
  wire       [3:0]    AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_robPtr;
  wire                AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_isFPR;
  wire                AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_hasException;
  wire       [7:0]    AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_exceptionCode;
  wire                AluIntEU_AluIntEuPlugin_setup_clearBusyPort_valid;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_setup_clearBusyPort_payload;
  wire                MulEU_MulEuPlugin_wakeupSourcePort_valid;
  wire       [5:0]    MulEU_MulEuPlugin_wakeupSourcePort_payload_physRegIdx;
  wire                MulEU_MulEuPlugin_gprReadPorts_0_valid;
  wire       [5:0]    MulEU_MulEuPlugin_gprReadPorts_0_address;
  wire       [31:0]   MulEU_MulEuPlugin_gprReadPorts_0_rsp;
  wire                MulEU_MulEuPlugin_gprReadPorts_1_valid;
  wire       [5:0]    MulEU_MulEuPlugin_gprReadPorts_1_address;
  wire       [31:0]   MulEU_MulEuPlugin_gprReadPorts_1_rsp;
  wire                MulEU_MulEuPlugin_gprWritePort_valid;
  wire       [5:0]    MulEU_MulEuPlugin_gprWritePort_address;
  wire       [31:0]   MulEU_MulEuPlugin_gprWritePort_data;
  wire                MulEU_MulEuPlugin_bypassOutputPort_valid;
  wire       [5:0]    MulEU_MulEuPlugin_bypassOutputPort_payload_physRegIdx;
  wire       [31:0]   MulEU_MulEuPlugin_bypassOutputPort_payload_physRegData;
  wire       [3:0]    MulEU_MulEuPlugin_bypassOutputPort_payload_robPtr;
  wire                MulEU_MulEuPlugin_bypassOutputPort_payload_isFPR;
  wire                MulEU_MulEuPlugin_bypassOutputPort_payload_hasException;
  wire       [7:0]    MulEU_MulEuPlugin_bypassOutputPort_payload_exceptionCode;
  wire                MulEU_MulEuPlugin_setup_clearBusyPort_valid;
  wire       [5:0]    MulEU_MulEuPlugin_setup_clearBusyPort_payload;
  wire                BranchEU_BranchEuPlugin_wakeupSourcePort_valid;
  wire       [5:0]    BranchEU_BranchEuPlugin_wakeupSourcePort_payload_physRegIdx;
  wire                BranchEU_BranchEuPlugin_gprReadPorts_0_valid;
  wire       [5:0]    BranchEU_BranchEuPlugin_gprReadPorts_0_address;
  wire       [31:0]   BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  wire                BranchEU_BranchEuPlugin_gprReadPorts_1_valid;
  wire       [5:0]    BranchEU_BranchEuPlugin_gprReadPorts_1_address;
  wire       [31:0]   BranchEU_BranchEuPlugin_gprReadPorts_1_rsp;
  wire                BranchEU_BranchEuPlugin_gprWritePort_valid;
  wire       [5:0]    BranchEU_BranchEuPlugin_gprWritePort_address;
  wire       [31:0]   BranchEU_BranchEuPlugin_gprWritePort_data;
  wire                BranchEU_BranchEuPlugin_bypassOutputPort_valid;
  wire       [5:0]    BranchEU_BranchEuPlugin_bypassOutputPort_payload_physRegIdx;
  wire       [31:0]   BranchEU_BranchEuPlugin_bypassOutputPort_payload_physRegData;
  wire       [3:0]    BranchEU_BranchEuPlugin_bypassOutputPort_payload_robPtr;
  wire                BranchEU_BranchEuPlugin_bypassOutputPort_payload_isFPR;
  wire                BranchEU_BranchEuPlugin_bypassOutputPort_payload_hasException;
  wire       [7:0]    BranchEU_BranchEuPlugin_bypassOutputPort_payload_exceptionCode;
  wire                BranchEU_BranchEuPlugin_setup_clearBusyPort_valid;
  wire       [5:0]    BranchEU_BranchEuPlugin_setup_clearBusyPort_payload;
  wire                LsuEU_LsuEuPlugin_wakeupSourcePort_valid;
  wire       [5:0]    LsuEU_LsuEuPlugin_wakeupSourcePort_payload_physRegIdx;
  wire                LsuEU_LsuEuPlugin_gprWritePort_valid;
  wire       [5:0]    LsuEU_LsuEuPlugin_gprWritePort_address;
  wire       [31:0]   LsuEU_LsuEuPlugin_gprWritePort_data;
  wire                LsuEU_LsuEuPlugin_bypassOutputPort_valid;
  wire       [5:0]    LsuEU_LsuEuPlugin_bypassOutputPort_payload_physRegIdx;
  wire       [31:0]   LsuEU_LsuEuPlugin_bypassOutputPort_payload_physRegData;
  wire       [3:0]    LsuEU_LsuEuPlugin_bypassOutputPort_payload_robPtr;
  wire                LsuEU_LsuEuPlugin_bypassOutputPort_payload_isFPR;
  wire                LsuEU_LsuEuPlugin_bypassOutputPort_payload_hasException;
  wire       [7:0]    LsuEU_LsuEuPlugin_bypassOutputPort_payload_exceptionCode;
  wire                LsuEU_LsuEuPlugin_setup_clearBusyPort_valid;
  wire       [5:0]    LsuEU_LsuEuPlugin_setup_clearBusyPort_payload;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_input_valid;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_input_ready;
  wire       [2:0]    LsuEU_LsuEuPlugin_hw_aguPort_input_payload_qPtr;
  wire       [5:0]    LsuEU_LsuEuPlugin_hw_aguPort_input_payload_basePhysReg;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_aguPort_input_payload_immediate;
  wire       [1:0]    LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_input_payload_usePc;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_aguPort_input_payload_pc;
  wire       [5:0]    LsuEU_LsuEuPlugin_hw_aguPort_input_payload_dataReg;
  wire       [3:0]    LsuEU_LsuEuPlugin_hw_aguPort_input_payload_robPtr;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isLoad;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isStore;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isFlush;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isIO;
  wire       [5:0]    LsuEU_LsuEuPlugin_hw_aguPort_input_payload_physDst;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_output_valid;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_output_ready;
  wire       [2:0]    LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException;
  wire       [1:0]    LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize;
  wire       [3:0]    LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask;
  wire       [5:0]    LsuEU_LsuEuPlugin_hw_aguPort_output_payload_basePhysReg;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc;
  wire       [3:0]    LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isStore;
  wire       [5:0]    LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_flush;
  wire                StoreBufferPlugin_hw_pushPortInst_valid;
  wire                StoreBufferPlugin_hw_pushPortInst_ready;
  wire       [31:0]   StoreBufferPlugin_hw_pushPortInst_payload_addr;
  wire       [31:0]   StoreBufferPlugin_hw_pushPortInst_payload_data;
  wire       [3:0]    StoreBufferPlugin_hw_pushPortInst_payload_be;
  wire       [3:0]    StoreBufferPlugin_hw_pushPortInst_payload_robPtr;
  wire       [1:0]    StoreBufferPlugin_hw_pushPortInst_payload_accessSize;
  wire                StoreBufferPlugin_hw_pushPortInst_payload_isFlush;
  wire                StoreBufferPlugin_hw_pushPortInst_payload_isIO;
  wire                StoreBufferPlugin_hw_pushPortInst_payload_hasEarlyException;
  wire       [7:0]    StoreBufferPlugin_hw_pushPortInst_payload_earlyExceptionCode;
  wire       [31:0]   StoreBufferPlugin_hw_bypassQueryAddrIn;
  wire       [1:0]    StoreBufferPlugin_hw_bypassQuerySizeIn;
  wire                StoreBufferPlugin_hw_bypassDataOutInst_valid;
  wire                StoreBufferPlugin_hw_bypassDataOutInst_payload_hit;
  wire       [31:0]   StoreBufferPlugin_hw_bypassDataOutInst_payload_data;
  wire       [3:0]    StoreBufferPlugin_hw_bypassDataOutInst_payload_hitMask;
  wire                StoreBufferPlugin_hw_sqQueryPort_cmd_valid;
  wire       [3:0]    StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr;
  wire       [31:0]   StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address;
  wire       [1:0]    StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size;
  wire                StoreBufferPlugin_hw_sqQueryPort_rsp_hit;
  wire       [31:0]   StoreBufferPlugin_hw_sqQueryPort_rsp_data;
  wire                StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreHasUnknownAddress;
  wire                StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreDataNotReady;
  wire                StoreBufferPlugin_hw_dCacheStorePort_cmd_valid;
  wire                StoreBufferPlugin_hw_dCacheStorePort_cmd_ready;
  reg        [31:0]   StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_address;
  reg        [31:0]   StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_data;
  reg        [3:0]    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_mask;
  reg                 StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_io;
  reg                 StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flush;
  reg                 StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flushFree;
  reg                 StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_prefetch;
  reg        [2:0]    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_id;
  wire                StoreBufferPlugin_hw_dCacheStorePort_rsp_valid;
  wire                StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_fault;
  wire                StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_redo;
  wire       [7:0]    StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_refillSlot;
  wire                StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_refillSlotAny;
  wire                StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_flush;
  wire                StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_prefetch;
  wire       [31:0]   StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_address;
  wire                StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_io;
  wire       [2:0]    StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_id;
  reg                 LoadQueuePlugin_hw_busyTableClearPort_valid;
  reg        [5:0]    LoadQueuePlugin_hw_busyTableClearPort_payload;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_cmd_valid;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_cmd_ready;
  wire       [31:0]   LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_virtual;
  wire       [1:0]    LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_redoOnDataHazard;
  wire       [2:0]    LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_transactionId;
  wire       [2:0]    LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_id;
  wire       [31:0]   LoadQueuePlugin_hw_dCacheLoadPort_translated_physical;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_translated_abord;
  wire       [2:0]    LoadQueuePlugin_hw_dCacheLoadPort_cancels;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_rsp_valid;
  wire       [31:0]   LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_data;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_fault;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_redo;
  wire       [7:0]    LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_refillSlot;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_refillSlotAny;
  wire       [2:0]    LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_id;
  reg                 LoadQueuePlugin_hw_prfWritePort_valid;
  reg        [5:0]    LoadQueuePlugin_hw_prfWritePort_address;
  reg        [31:0]   LoadQueuePlugin_hw_prfWritePort_data;
  reg                 LoadQueuePlugin_hw_wakeupPort_valid;
  reg        [5:0]    LoadQueuePlugin_hw_wakeupPort_payload_physRegIdx;
  wire                _zz_LoadQueuePlugin_logic_loadQueue_mmioCmdFired;
  reg                 CheckpointManagerPlugin_setup_btRestorePort_valid;
  reg        [63:0]   CheckpointManagerPlugin_setup_btRestorePort_payload_busyBits;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid;
  wire       [5:0]    LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_address;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp;
  wire                LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_valid;
  wire       [5:0]    LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_address;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp;
  wire                LsuEU_LsuEuPlugin_hw_lqPushPort_valid;
  wire                LsuEU_LsuEuPlugin_hw_lqPushPort_ready;
  wire       [3:0]    LsuEU_LsuEuPlugin_hw_lqPushPort_payload_robPtr;
  wire       [5:0]    LsuEU_LsuEuPlugin_hw_lqPushPort_payload_pdest;
  wire       [31:0]   LsuEU_LsuEuPlugin_hw_lqPushPort_payload_address;
  wire                LsuEU_LsuEuPlugin_hw_lqPushPort_payload_isIO;
  wire       [1:0]    LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size;
  wire                LsuEU_LsuEuPlugin_hw_lqPushPort_payload_hasEarlyException;
  wire       [7:0]    LsuEU_LsuEuPlugin_hw_lqPushPort_payload_earlyExceptionCode;
  wire                LinkerPlugin_logic_allWakeupFlows_0_valid;
  wire       [5:0]    LinkerPlugin_logic_allWakeupFlows_0_payload_physRegIdx;
  wire                LinkerPlugin_logic_allWakeupFlows_1_valid;
  wire       [5:0]    LinkerPlugin_logic_allWakeupFlows_1_payload_physRegIdx;
  wire                LinkerPlugin_logic_allWakeupFlows_2_valid;
  wire       [5:0]    LinkerPlugin_logic_allWakeupFlows_2_payload_physRegIdx;
  wire                LinkerPlugin_logic_allWakeupFlows_3_valid;
  wire       [5:0]    LinkerPlugin_logic_allWakeupFlows_3_payload_physRegIdx;
  wire                LinkerPlugin_logic_allWakeupFlows_4_valid;
  wire       [5:0]    LinkerPlugin_logic_allWakeupFlows_4_payload_physRegIdx;
  wire                AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_valid;
  wire                AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_ready;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_physRegIdx;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_physRegData;
  wire       [3:0]    AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_robPtr;
  wire                AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_isFPR;
  wire                AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_hasException;
  wire       [7:0]    AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_exceptionCode;
  wire                MulEU_MulEuPlugin_bypassOutputPort_toStream_valid;
  wire                MulEU_MulEuPlugin_bypassOutputPort_toStream_ready;
  wire       [5:0]    MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_physRegIdx;
  wire       [31:0]   MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_physRegData;
  wire       [3:0]    MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_robPtr;
  wire                MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_isFPR;
  wire                MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_hasException;
  wire       [7:0]    MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_exceptionCode;
  wire                BranchEU_BranchEuPlugin_bypassOutputPort_toStream_valid;
  wire                BranchEU_BranchEuPlugin_bypassOutputPort_toStream_ready;
  wire       [5:0]    BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_physRegIdx;
  wire       [31:0]   BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_physRegData;
  wire       [3:0]    BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_robPtr;
  wire                BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_isFPR;
  wire                BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_hasException;
  wire       [7:0]    BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_exceptionCode;
  wire                io_output_combStage_valid;
  wire                io_output_combStage_ready;
  wire       [5:0]    io_output_combStage_payload_physRegIdx;
  wire       [31:0]   io_output_combStage_payload_physRegData;
  wire       [3:0]    io_output_combStage_payload_robPtr;
  wire                io_output_combStage_payload_isFPR;
  wire                io_output_combStage_payload_hasException;
  wire       [7:0]    io_output_combStage_payload_exceptionCode;
  wire                AguPlugin_logic_bypassFlow_valid;
  wire       [5:0]    AguPlugin_logic_bypassFlow_payload_physRegIdx;
  wire       [31:0]   AguPlugin_logic_bypassFlow_payload_physRegData;
  wire       [3:0]    AguPlugin_logic_bypassFlow_payload_robPtr;
  wire                AguPlugin_logic_bypassFlow_payload_isFPR;
  wire                AguPlugin_logic_bypassFlow_payload_hasException;
  wire       [7:0]    AguPlugin_logic_bypassFlow_payload_exceptionCode;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_0;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_1;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_2;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_3;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_4;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_5;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_6;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_7;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_8;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_9;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_10;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_11;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_12;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_13;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_14;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_15;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_16;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_17;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_18;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_19;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_20;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_21;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_22;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_23;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_24;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_25;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_26;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_27;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_28;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_29;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_30;
  reg        [5:0]    CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_31;
  reg        [63:0]   CheckpointManagerPlugin_logic_storedBtCheckpoint_busyBits;
  reg                 CheckpointManagerPlugin_logic_hasValidCheckpoint;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_0;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_1;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_2;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_3;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_4;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_5;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_6;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_7;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_8;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_9;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_10;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_11;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_12;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_13;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_14;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_15;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_16;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_17;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_18;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_19;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_20;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_21;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_22;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_23;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_24;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_25;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_26;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_27;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_28;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_29;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_30;
  wire       [5:0]    CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_31;
  reg        [63:0]   CheckpointManagerPlugin_logic_initialFreeMask;
  wire       [63:0]   CheckpointManagerPlugin_logic_initialBtCheckpoint_busyBits;
  wire                CommitPlugin_logic_s0_isMispredictedBranch;
  reg                 CommitPlugin_logic_s0_commitAckMasks_0;
  wire                when_CommitPlugin_l203;
  wire                when_CommitPlugin_l216;
  wire                when_CommitPlugin_l227;
  wire                when_CommitPlugin_l265;
  wire       [0:0]    CommitPlugin_logic_s0_committedThisCycle_comb;
  wire       [0:0]    CommitPlugin_logic_s0_recycledThisCycle_comb;
  wire       [0:0]    CommitPlugin_logic_s0_flushedThisCycle_comb;
  wire       [31:0]   CommitPlugin_logic_s0_commitPcs_0;
  wire       [31:0]   CommitPlugin_logic_s0_maxCommitPcThisCycle;
  wire                CommitPlugin_logic_s0_anyCommitOOB;
  wire                CommitPlugin_logic_s0_commitSlotLogs_0_valid;
  wire                CommitPlugin_logic_s0_commitSlotLogs_0_canCommit;
  wire                CommitPlugin_logic_s0_commitSlotLogs_0_doCommit;
  wire       [3:0]    CommitPlugin_logic_s0_commitSlotLogs_0_robPtr;
  wire       [5:0]    CommitPlugin_logic_s0_commitSlotLogs_0_oldPhysDest;
  wire                CommitPlugin_logic_s0_commitSlotLogs_0_allocatesPhysDest;
  reg        [0:0]    CommitPlugin_logic_s1_s1_committedThisCycle;
  reg        [0:0]    CommitPlugin_logic_s1_s1_recycledThisCycle;
  reg        [0:0]    CommitPlugin_logic_s1_s1_flushedThisCycle;
  reg        [31:0]   CommitPlugin_logic_s1_s1_maxCommitPcThisCycle;
  reg                 CommitPlugin_logic_s1_s1_anyCommitOOB;
  wire                CommitPlugin_logic_s1_s1_hasCommitsThisCycle;
  wire                when_CommitPlugin_l317;
  wire       [4:0]    _zz_when_Debug_l71_6;
  wire                when_Debug_l71_5;
  wire       [7:0]    _zz_26;
  reg        [31:0]   CommitPlugin_logic_counter;
  wire       [31:0]   DecodePlugin_logic_decodedUopsOutputVec_0_pc;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_isValid;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_uopCode;
  wire       [3:0]    DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_isa;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_archDest_idx;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_writeArchDestEn;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_idx;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_useArchSrc1;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_idx;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_useArchSrc2;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_usePcForAddr;
  wire       [31:0]   DecodePlugin_logic_decodedUopsOutputVec_0_imm;
  wire       [2:0]    DecodePlugin_logic_decodedUopsOutputVec_0_immUsage;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_valid;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isSub;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isAdd;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isSigned;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_valid;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isRight;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isArithmetic;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isRotate;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isDoubleWord;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_valid;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isDiv;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isSigned;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isWordOp;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isSignedLoad;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isStore;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isLoadLinked;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isStoreCond;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_atomicOp;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isFence;
  wire       [7:0]    DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_fenceMode;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isCacheOp;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_cacheOpType;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isPrefetch;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isJump;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isLink;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_idx;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isIndirect;
  wire       [2:0]    DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_laCfIdx;
  wire       [3:0]    DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_opType;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest;
  wire       [2:0]    DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_roundingMode;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_isIntegerDest;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_isSignedCvt;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fcmpCond;
  wire       [13:0]   DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_csrAddr;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isWrite;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isRead;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isExchange;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_useUimmAsSrc;
  wire       [19:0]   DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_sysCode;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_isExceptionReturn;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_isTlbOp;
  wire       [3:0]    DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_tlbOpType;
  wire       [1:0]    DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_hasDecodeException;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_isMicrocode;
  wire       [7:0]    DecodePlugin_logic_decodedUopsOutputVec_0_microcodeEntry;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_isSerializing;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_isBranchOrJump;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken;
  wire       [31:0]   DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target;
  wire                DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted;
  reg                 _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isValid;
  reg        [4:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode;
  wire       [3:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype;
  wire                _zz_DecodePlugin_logic_decodedUopsOutputVec_0_writeArchDestEn;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype;
  wire       [4:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_idx;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype;
  wire       [2:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size;
  wire       [4:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest;
  reg        [1:0]    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode;
  reg                 _zz_DecodePlugin_logic_decodedUopsOutputVec_0_hasDecodeException;
  reg                 _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken;
  reg        [31:0]   _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target;
  reg                 _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [4:0]    DecodePlugin_logic_debugLA32RDecodedPhysSrc2_idx;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [1:0]    DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [31:0]   DecodePlugin_logic_debugLA32RRawInstruction;
  wire                when_DecodePlugin_l66;
  wire                when_DecodePlugin_l79;
  wire                when_DecodePlugin_l85;
  wire                when_DecodePlugin_l117;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                RenamePlugin_logic_s2_logic_allocationOk;
  wire                when_RenamePlugin_l83;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                s2_RobAlloc_haltRequest_RenamePlugin_l85;
  wire                s2_RobAlloc_haltRequest_RobAllocPlugin_l30;
  wire       [31:0]   RobAllocPlugin_logic_allocatedUops_0_decoded_pc;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_isValid;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode;
  wire       [3:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_isa;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_idx;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_writeArchDestEn;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_idx;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_useArchSrc1;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_idx;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_useArchSrc2;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_usePcForAddr;
  wire       [31:0]   RobAllocPlugin_logic_allocatedUops_0_decoded_imm;
  wire       [2:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_valid;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isSub;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isAdd;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isSigned;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_valid;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isRight;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isArithmetic;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isRotate;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isDoubleWord;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_valid;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isDiv;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isSigned;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isWordOp;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isSignedLoad;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isStore;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isLoadLinked;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isStoreCond;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_atomicOp;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isFence;
  wire       [7:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_fenceMode;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isCacheOp;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_cacheOpType;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isPrefetch;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isJump;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isLink;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isIndirect;
  wire       [2:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_laCfIdx;
  wire       [3:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_opType;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest;
  wire       [2:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_roundingMode;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_isIntegerDest;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_isSignedCvt;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fcmpCond;
  wire       [13:0]   RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_csrAddr;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isWrite;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isRead;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isExchange;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_useUimmAsSrc;
  wire       [19:0]   RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_sysCode;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_isExceptionReturn;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_isTlbOp;
  wire       [3:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_tlbOpType;
  wire       [1:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_hasDecodeException;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_isMicrocode;
  wire       [7:0]    RobAllocPlugin_logic_allocatedUops_0_decoded_microcodeEntry;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_isSerializing;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_isBranchOrJump;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_isTaken;
  wire       [31:0]   RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_target;
  wire                RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_wasPredicted;
  wire       [5:0]    RobAllocPlugin_logic_allocatedUops_0_rename_physSrc1_idx;
  wire                RobAllocPlugin_logic_allocatedUops_0_rename_physSrc1IsFpr;
  wire       [5:0]    RobAllocPlugin_logic_allocatedUops_0_rename_physSrc2_idx;
  wire                RobAllocPlugin_logic_allocatedUops_0_rename_physSrc2IsFpr;
  wire       [5:0]    RobAllocPlugin_logic_allocatedUops_0_rename_physDest_idx;
  wire                RobAllocPlugin_logic_allocatedUops_0_rename_physDestIsFpr;
  wire       [5:0]    RobAllocPlugin_logic_allocatedUops_0_rename_oldPhysDest_idx;
  wire                RobAllocPlugin_logic_allocatedUops_0_rename_oldPhysDestIsFpr;
  wire                RobAllocPlugin_logic_allocatedUops_0_rename_allocatesPhysDest;
  wire                RobAllocPlugin_logic_allocatedUops_0_rename_writesToPhysReg;
  wire       [3:0]    RobAllocPlugin_logic_allocatedUops_0_robPtr;
  wire       [15:0]   RobAllocPlugin_logic_allocatedUops_0_uniqueId;
  wire                RobAllocPlugin_logic_allocatedUops_0_dispatched;
  wire                RobAllocPlugin_logic_allocatedUops_0_executed;
  wire                RobAllocPlugin_logic_allocatedUops_0_hasException;
  wire       [7:0]    RobAllocPlugin_logic_allocatedUops_0_exceptionCode;
  wire                DispatchPlugin_logic_iqRegs_0_1_valid;
  wire                DispatchPlugin_logic_iqRegs_0_1_ready;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_pc;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isValid;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_writeArchDestEn;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_useArchSrc1;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_useArchSrc2;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_usePcForAddr;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_imm;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isSub;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isAdd;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isRight;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isArithmetic;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isRotate;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isDiv;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isSigned;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isSignedLoad;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isStore;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isLoadLinked;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_atomicOp;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isFence;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_fenceMode;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_cacheOpType;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isJump;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_roundingMode;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_csrAddr;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isWrite;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isRead;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isExchange;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_sysCode;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_hasDecodeException;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isMicrocode;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_microcodeEntry;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isSerializing;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isBranchOrJump;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_target;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc1_idx;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc1IsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc2_idx;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc2IsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physDest_idx;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physDestIsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_oldPhysDest_idx;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_oldPhysDestIsFpr;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_allocatesPhysDest;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_writesToPhysReg;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_robPtr;
  reg        [15:0]   DispatchPlugin_logic_iqRegs_0_1_payload_uop_uniqueId;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_dispatched;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_executed;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_uop_hasException;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_0_1_payload_uop_exceptionCode;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_src1InitialReady;
  reg                 DispatchPlugin_logic_iqRegs_0_1_payload_src2InitialReady;
  wire                DispatchPlugin_logic_iqRegs_1_1_valid;
  wire                DispatchPlugin_logic_iqRegs_1_1_ready;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_pc;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isValid;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_writeArchDestEn;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_useArchSrc1;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_useArchSrc2;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_usePcForAddr;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_imm;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isSub;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isAdd;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isRight;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isArithmetic;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isRotate;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isDiv;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isSigned;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isSignedLoad;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isStore;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isLoadLinked;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_atomicOp;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isFence;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_fenceMode;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_cacheOpType;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isJump;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_roundingMode;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_csrAddr;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isWrite;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isRead;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isExchange;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_sysCode;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_hasDecodeException;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isMicrocode;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_microcodeEntry;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isSerializing;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isBranchOrJump;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_target;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc1_idx;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc1IsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc2_idx;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc2IsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physDest_idx;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physDestIsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_oldPhysDest_idx;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_oldPhysDestIsFpr;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_allocatesPhysDest;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_writesToPhysReg;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_robPtr;
  reg        [15:0]   DispatchPlugin_logic_iqRegs_1_1_payload_uop_uniqueId;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_dispatched;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_executed;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_uop_hasException;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_1_1_payload_uop_exceptionCode;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_src1InitialReady;
  reg                 DispatchPlugin_logic_iqRegs_1_1_payload_src2InitialReady;
  wire                DispatchPlugin_logic_iqRegs_2_1_valid;
  wire                DispatchPlugin_logic_iqRegs_2_1_ready;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_pc;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isValid;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_writeArchDestEn;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_useArchSrc1;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_useArchSrc2;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_usePcForAddr;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_imm;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isSub;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isAdd;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isRight;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isArithmetic;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isRotate;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isDiv;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isSigned;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isSignedLoad;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isStore;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isLoadLinked;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_atomicOp;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isFence;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_fenceMode;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_cacheOpType;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isJump;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_roundingMode;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_csrAddr;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isWrite;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isRead;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isExchange;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_sysCode;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_hasDecodeException;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isMicrocode;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_microcodeEntry;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isSerializing;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isBranchOrJump;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_target;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc1_idx;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc1IsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc2_idx;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc2IsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physDest_idx;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physDestIsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_oldPhysDest_idx;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_oldPhysDestIsFpr;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_allocatesPhysDest;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_writesToPhysReg;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_robPtr;
  reg        [15:0]   DispatchPlugin_logic_iqRegs_2_1_payload_uop_uniqueId;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_dispatched;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_executed;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_uop_hasException;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_2_1_payload_uop_exceptionCode;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_src1InitialReady;
  reg                 DispatchPlugin_logic_iqRegs_2_1_payload_src2InitialReady;
  wire                DispatchPlugin_logic_iqRegs_3_1_valid;
  wire                DispatchPlugin_logic_iqRegs_3_1_ready;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_pc;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isValid;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_writeArchDestEn;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_useArchSrc1;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_useArchSrc2;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_usePcForAddr;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_imm;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isSub;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isAdd;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isRight;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isArithmetic;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isRotate;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_valid;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isDiv;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isSigned;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isSignedLoad;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isStore;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isLoadLinked;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_atomicOp;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isFence;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_fenceMode;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_cacheOpType;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isJump;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_roundingMode;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_csrAddr;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isWrite;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isRead;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isExchange;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_sysCode;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_hasDecodeException;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isMicrocode;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_microcodeEntry;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isSerializing;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isBranchOrJump;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_target;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc1_idx;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc1IsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc2_idx;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc2IsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physDest_idx;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physDestIsFpr;
  reg        [5:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_oldPhysDest_idx;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_oldPhysDestIsFpr;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_allocatesPhysDest;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_writesToPhysReg;
  reg        [3:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_robPtr;
  reg        [15:0]   DispatchPlugin_logic_iqRegs_3_1_payload_uop_uniqueId;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_dispatched;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_executed;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_uop_hasException;
  reg        [7:0]    DispatchPlugin_logic_iqRegs_3_1_payload_uop_exceptionCode;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_src1InitialReady;
  reg                 DispatchPlugin_logic_iqRegs_3_1_payload_src2InitialReady;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_valid;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_ready;
  wire       [3:0]    AluIntEU_AluIntEuPlugin_euInputPort_payload_robPtr;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_euInputPort_payload_physDest_idx;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_physDestIsFpr;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_writesToPhysReg;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_useSrc1;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Data;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Tag;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Ready;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_src1IsFpr;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_useSrc2;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Data;
  wire       [5:0]    AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Tag;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Ready;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_src2IsFpr;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_valid;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isSub;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isAdd;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isSigned;
  wire       [1:0]    AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_valid;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isRight;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isArithmetic;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isRotate;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isDoubleWord;
  wire       [31:0]   AluIntEU_AluIntEuPlugin_euInputPort_payload_imm;
  wire       [2:0]    AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage;
  wire                AluIntEU_AluIntEuPlugin_euInputPort_fire;
  wire                MulEU_MulEuPlugin_euInputPort_valid;
  wire                MulEU_MulEuPlugin_euInputPort_ready;
  wire       [31:0]   MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_pc;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isValid;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode;
  wire       [3:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_idx;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_writeArchDestEn;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_idx;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_useArchSrc1;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_idx;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_useArchSrc2;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_usePcForAddr;
  wire       [31:0]   MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_imm;
  wire       [2:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_valid;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_isSub;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_isAdd;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_isSigned;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_valid;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_isRight;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_isArithmetic;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_isRotate;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_isDoubleWord;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_mulDivCtrl_valid;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_mulDivCtrl_isDiv;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_mulDivCtrl_isSigned;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_mulDivCtrl_isWordOp;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isSignedLoad;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isStore;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isLoadLinked;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isStoreCond;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_atomicOp;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isFence;
  wire       [7:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_fenceMode;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isCacheOp;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_cacheOpType;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isPrefetch;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_isJump;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_isLink;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_isIndirect;
  wire       [2:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_laCfIdx;
  wire       [3:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_opType;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest;
  wire       [2:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_roundingMode;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_isIntegerDest;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_isSignedCvt;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  wire       [4:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fcmpCond;
  wire       [13:0]   MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_csrAddr;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_isWrite;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_isRead;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_isExchange;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  wire       [19:0]   MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_sysCtrl_sysCode;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_sysCtrl_isExceptionReturn;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_sysCtrl_isTlbOp;
  wire       [3:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_sysCtrl_tlbOpType;
  wire       [1:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_hasDecodeException;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isMicrocode;
  wire       [7:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_microcodeEntry;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isSerializing;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isBranchOrJump;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchPrediction_isTaken;
  wire       [31:0]   MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchPrediction_target;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchPrediction_wasPredicted;
  wire       [5:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physSrc1_idx;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physSrc1IsFpr;
  wire       [5:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physSrc2_idx;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physSrc2IsFpr;
  wire       [5:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physDest_idx;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physDestIsFpr;
  wire       [5:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_rename_oldPhysDest_idx;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_rename_oldPhysDestIsFpr;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_rename_allocatesPhysDest;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_rename_writesToPhysReg;
  wire       [3:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_robPtr;
  wire       [15:0]   MulEU_MulEuPlugin_euInputPort_payload_uop_uniqueId;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_dispatched;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_executed;
  wire                MulEU_MulEuPlugin_euInputPort_payload_uop_hasException;
  wire       [7:0]    MulEU_MulEuPlugin_euInputPort_payload_uop_exceptionCode;
  wire       [3:0]    MulEU_MulEuPlugin_euInputPort_payload_robPtr;
  wire       [5:0]    MulEU_MulEuPlugin_euInputPort_payload_physDest_idx;
  wire                MulEU_MulEuPlugin_euInputPort_payload_physDestIsFpr;
  wire                MulEU_MulEuPlugin_euInputPort_payload_writesToPhysReg;
  wire                MulEU_MulEuPlugin_euInputPort_payload_useSrc1;
  wire       [31:0]   MulEU_MulEuPlugin_euInputPort_payload_src1Data;
  wire       [5:0]    MulEU_MulEuPlugin_euInputPort_payload_src1Tag;
  wire                MulEU_MulEuPlugin_euInputPort_payload_src1Ready;
  wire                MulEU_MulEuPlugin_euInputPort_payload_src1IsFpr;
  wire                MulEU_MulEuPlugin_euInputPort_payload_useSrc2;
  wire       [31:0]   MulEU_MulEuPlugin_euInputPort_payload_src2Data;
  wire       [5:0]    MulEU_MulEuPlugin_euInputPort_payload_src2Tag;
  wire                MulEU_MulEuPlugin_euInputPort_payload_src2Ready;
  wire                MulEU_MulEuPlugin_euInputPort_payload_src2IsFpr;
  wire                MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_valid;
  wire                MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isDiv;
  wire                MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isSigned;
  wire                MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isWordOp;
  wire                MulEU_MulEuPlugin_euInputPort_fire;
  wire                BranchEU_BranchEuPlugin_euInputPort_valid;
  wire                BranchEU_BranchEuPlugin_euInputPort_ready;
  wire       [3:0]    BranchEU_BranchEuPlugin_euInputPort_payload_robPtr;
  wire       [5:0]    BranchEU_BranchEuPlugin_euInputPort_payload_physDest_idx;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_physDestIsFpr;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_writesToPhysReg;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_useSrc1;
  wire       [31:0]   BranchEU_BranchEuPlugin_euInputPort_payload_src1Data;
  wire       [5:0]    BranchEU_BranchEuPlugin_euInputPort_payload_src1Tag;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_src1Ready;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_src1IsFpr;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_useSrc2;
  wire       [31:0]   BranchEU_BranchEuPlugin_euInputPort_payload_src2Data;
  wire       [5:0]    BranchEU_BranchEuPlugin_euInputPort_payload_src2Tag;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_src2Ready;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_src2IsFpr;
  wire       [4:0]    BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isJump;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isLink;
  wire       [4:0]    BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_idx;
  wire       [1:0]    BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isIndirect;
  wire       [2:0]    BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_laCfIdx;
  wire       [31:0]   BranchEU_BranchEuPlugin_euInputPort_payload_imm;
  wire       [31:0]   BranchEU_BranchEuPlugin_euInputPort_payload_pc;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_isTaken;
  wire       [31:0]   BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_target;
  wire                BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_wasPredicted;
  wire                BranchEU_BranchEuPlugin_euInputPort_fire;
  wire                LsuEU_LsuEuPlugin_euInputPort_valid;
  wire                LsuEU_LsuEuPlugin_euInputPort_ready;
  wire       [3:0]    LsuEU_LsuEuPlugin_euInputPort_payload_robPtr;
  wire       [5:0]    LsuEU_LsuEuPlugin_euInputPort_payload_physDest_idx;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_physDestIsFpr;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_writesToPhysReg;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_useSrc1;
  wire       [31:0]   LsuEU_LsuEuPlugin_euInputPort_payload_src1Data;
  wire       [5:0]    LsuEU_LsuEuPlugin_euInputPort_payload_src1Tag;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_src1Ready;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_src1IsFpr;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_useSrc2;
  wire       [31:0]   LsuEU_LsuEuPlugin_euInputPort_payload_src2Data;
  wire       [5:0]    LsuEU_LsuEuPlugin_euInputPort_payload_src2Tag;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_src2Ready;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_src2IsFpr;
  wire       [1:0]    LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isSignedLoad;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isStore;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isLoadLinked;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isStoreCond;
  wire       [4:0]    LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_atomicOp;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isFence;
  wire       [7:0]    LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_fenceMode;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isCacheOp;
  wire       [4:0]    LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_cacheOpType;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isPrefetch;
  wire       [31:0]   LsuEU_LsuEuPlugin_euInputPort_payload_imm;
  wire                LsuEU_LsuEuPlugin_euInputPort_payload_usePc;
  wire       [31:0]   LsuEU_LsuEuPlugin_euInputPort_payload_pcData;
  wire                LsuEU_LsuEuPlugin_euInputPort_fire;
  wire       [4:0]    _zz_when_Debug_l71_7;
  wire                when_Debug_l71_6;
  wire                DispatchPlugin_logic_physSrc1ConflictS1;
  wire                DispatchPlugin_logic_physSrc1ConflictS2;
  wire                DispatchPlugin_logic_physSrc2ConflictS1;
  wire                DispatchPlugin_logic_physSrc2ConflictS2;
  wire                DispatchPlugin_logic_src1SetBypass;
  wire                DispatchPlugin_logic_src2SetBypass;
  wire                DispatchPlugin_logic_src1ReadyCandidate;
  wire                DispatchPlugin_logic_src1InitialReady;
  wire                DispatchPlugin_logic_src2ReadyCandidate;
  wire                DispatchPlugin_logic_src2InitialReady;
  wire       [3:0]    DispatchPlugin_logic_dispatchOH;
  wire                _zz_DispatchPlugin_logic_destinationIqReady;
  wire                _zz_DispatchPlugin_logic_destinationIqReady_1;
  wire                _zz_DispatchPlugin_logic_destinationIqReady_2;
  wire                DispatchPlugin_logic_destinationIqReady;
  wire                s3_Dispatch_haltRequest_DispatchPlugin_l78;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    DispatchPlugin_logic_debugDispatchedUopSrc2_iq0;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    DispatchPlugin_logic_debugDispatchedUopSrc1_iq0;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    DispatchPlugin_logic_debugDispatchedUopSrc2_iq1;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    DispatchPlugin_logic_debugDispatchedUopSrc1_iq1;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    DispatchPlugin_logic_debugDispatchedUopSrc2_iq2;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    DispatchPlugin_logic_debugDispatchedUopSrc1_iq2;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    DispatchPlugin_logic_debugDispatchedUopSrc2_iq3;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    DispatchPlugin_logic_debugDispatchedUopSrc1_iq3;
  wire                when_DispatchPlugin_l100;
  wire       [31:0]   CoreNSCSCCSetupPlugin_logic_instructionVec_0;
  wire       [31:0]   CoreNSCSCCSetupPlugin_logic_instructionVec_1;
  wire       [31:0]   CoreNSCSCCSetupPlugin_logic_instructionVec_2;
  wire       [31:0]   CoreNSCSCCSetupPlugin_logic_instructionVec_3;
  reg                 DebugDisplayPlugin_logic_displayArea_dpToggle;
  wire                s0_Dispatch_valid;
  reg                 _zz_s1_ReadRegs_valid;
  reg                 s1_ReadRegs_valid;
  reg                 _zz_s2_Execute_valid;
  reg                 s2_Execute_valid;
  reg                 _zz_s3_Writeback_valid;
  reg                 s3_Writeback_valid;
  wire                s1_ReadRegs_isFiring;
  wire       [31:0]   _zz_io_iqEntryIn_payload_src2Data_1;
  wire                s2_Execute_isFiring;
  wire       [2:0]    _zz_51;
  wire                s3_Writeback_isFiring;
  wire                when_Connection_l66_1;
  wire                when_Connection_l66_2;
  wire                when_EuBasePlugin_l230;
  wire                AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes;
  wire                AluIntEU_AluIntEuPlugin_logicPhase_completesSuccessfully;
  wire       [4:0]    _zz_when_Debug_l71_8;
  wire                when_Debug_l71_7;
  wire                when_EuBasePlugin_l300;
  wire                mul_s0_Dispatch_valid;
  reg                 _zz_mul_s1_ReadRegs_valid;
  reg                 mul_s1_ReadRegs_valid;
  reg                 _zz_mul_s2_Execute_valid;
  reg                 mul_s2_Execute_valid;
  reg                 _zz_mul_s3_Execute_valid;
  reg                 mul_s3_Execute_valid;
  reg                 _zz_mul_s4_Execute_valid;
  reg                 mul_s4_Execute_valid;
  reg                 _zz_mul_s5_Execute_valid;
  reg                 mul_s5_Execute_valid;
  reg                 _zz_mul_s6_Execute_valid;
  reg                 mul_s6_Execute_valid;
  reg                 _zz_mul_s7_Writeback_valid;
  reg                 mul_s7_Writeback_valid;
  wire                mul_s1_ReadRegs_isFiring;
  wire                mul_s2_Execute_isFiring;
  wire                mul_s7_Writeback_isFiring;
  wire                when_Connection_l66_3;
  wire                when_Connection_l66_4;
  wire                when_Connection_l66_5;
  wire                when_Connection_l66_6;
  wire                when_Connection_l66_7;
  wire                when_Connection_l66_8;
  wire                when_EuBasePlugin_l230_1;
  wire                MulEU_MulEuPlugin_logicPhase_executionCompletes;
  wire                MulEU_MulEuPlugin_logicPhase_completesSuccessfully;
  wire       [4:0]    _zz_when_Debug_l71_9;
  wire                when_Debug_l71_8;
  wire                when_EuBasePlugin_l300_1;
  wire                s0_Dispatch_valid_1;
  reg                 _zz_s1_Calc_valid;
  reg                 s1_Calc_valid;
  reg                 _zz_s2_Select_valid;
  reg                 s2_Select_valid;
  reg                 _zz_s3_Result_valid;
  reg                 s3_Result_valid;
  wire                s0_Dispatch_isFiring;
  wire                s1_Calc_isFiring;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_data_3;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_data_4;
  wire       [1:0]    switch_BranchEuPlugin_l133;
  wire                s2_Select_isFiring;
  wire       [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_data_5;
  reg        [31:0]   _zz_BranchEU_BranchEuPlugin_euResult_data_6;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_isTaken_1;
  reg                 _zz_BranchEU_BranchEuPlugin_euResult_isMispredictedBranch_1;
  wire                _zz_52;
  wire                s3_Result_isFiring;
  wire                when_Connection_l66_9;
  wire                when_Connection_l66_10;
  wire                when_EuBasePlugin_l230_2;
  wire                BranchEU_BranchEuPlugin_logicPhase_executionCompletes;
  wire                BranchEU_BranchEuPlugin_logicPhase_completesSuccessfully;
  wire       [4:0]    _zz_when_Debug_l71_10;
  wire                when_Debug_l71_9;
  wire                when_EuBasePlugin_l300_2;
  wire       [1:0]    _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize;
  wire                LsuEU_LsuEuPlugin_euInputPort_translated_valid;
  wire                LsuEU_LsuEuPlugin_euInputPort_translated_ready;
  wire       [2:0]    LsuEU_LsuEuPlugin_euInputPort_translated_payload_qPtr;
  wire       [5:0]    LsuEU_LsuEuPlugin_euInputPort_translated_payload_basePhysReg;
  wire       [31:0]   LsuEU_LsuEuPlugin_euInputPort_translated_payload_immediate;
  wire       [1:0]    LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize;
  wire                LsuEU_LsuEuPlugin_euInputPort_translated_payload_usePc;
  wire       [31:0]   LsuEU_LsuEuPlugin_euInputPort_translated_payload_pc;
  wire       [5:0]    LsuEU_LsuEuPlugin_euInputPort_translated_payload_dataReg;
  wire       [3:0]    LsuEU_LsuEuPlugin_euInputPort_translated_payload_robPtr;
  wire                LsuEU_LsuEuPlugin_euInputPort_translated_payload_isLoad;
  wire                LsuEU_LsuEuPlugin_euInputPort_translated_payload_isStore;
  wire                LsuEU_LsuEuPlugin_euInputPort_translated_payload_isFlush;
  wire                LsuEU_LsuEuPlugin_euInputPort_translated_payload_isIO;
  wire       [5:0]    LsuEU_LsuEuPlugin_euInputPort_translated_payload_physDst;
  wire                io_outputs_0_combStage_valid;
  wire                io_outputs_0_combStage_ready;
  wire       [2:0]    io_outputs_0_combStage_payload_qPtr;
  wire       [31:0]   io_outputs_0_combStage_payload_address;
  wire                io_outputs_0_combStage_payload_alignException;
  wire       [1:0]    io_outputs_0_combStage_payload_accessSize;
  wire       [3:0]    io_outputs_0_combStage_payload_storeMask;
  wire       [5:0]    io_outputs_0_combStage_payload_basePhysReg;
  wire       [31:0]   io_outputs_0_combStage_payload_immediate;
  wire                io_outputs_0_combStage_payload_usePc;
  wire       [31:0]   io_outputs_0_combStage_payload_pc;
  wire       [3:0]    io_outputs_0_combStage_payload_robPtr;
  wire                io_outputs_0_combStage_payload_isLoad;
  wire                io_outputs_0_combStage_payload_isStore;
  wire       [5:0]    io_outputs_0_combStage_payload_physDst;
  wire       [31:0]   io_outputs_0_combStage_payload_storeData;
  wire                io_outputs_0_combStage_payload_isFlush;
  wire                io_outputs_0_combStage_payload_isIO;
  wire                io_outputs_1_combStage_valid;
  wire                io_outputs_1_combStage_ready;
  wire       [2:0]    io_outputs_1_combStage_payload_qPtr;
  wire       [31:0]   io_outputs_1_combStage_payload_address;
  wire                io_outputs_1_combStage_payload_alignException;
  wire       [1:0]    io_outputs_1_combStage_payload_accessSize;
  wire       [3:0]    io_outputs_1_combStage_payload_storeMask;
  wire       [5:0]    io_outputs_1_combStage_payload_basePhysReg;
  wire       [31:0]   io_outputs_1_combStage_payload_immediate;
  wire                io_outputs_1_combStage_payload_usePc;
  wire       [31:0]   io_outputs_1_combStage_payload_pc;
  wire       [3:0]    io_outputs_1_combStage_payload_robPtr;
  wire                io_outputs_1_combStage_payload_isLoad;
  wire                io_outputs_1_combStage_payload_isStore;
  wire       [5:0]    io_outputs_1_combStage_payload_physDst;
  wire       [31:0]   io_outputs_1_combStage_payload_storeData;
  wire                io_outputs_1_combStage_payload_isFlush;
  wire                io_outputs_1_combStage_payload_isIO;
  wire       [1:0]    _zz_io_outputs_0_combStage_translated_payload_size;
  wire                io_outputs_0_combStage_translated_valid;
  wire                io_outputs_0_combStage_translated_ready;
  wire       [3:0]    io_outputs_0_combStage_translated_payload_robPtr;
  wire       [5:0]    io_outputs_0_combStage_translated_payload_pdest;
  wire       [31:0]   io_outputs_0_combStage_translated_payload_address;
  wire                io_outputs_0_combStage_translated_payload_isIO;
  wire       [1:0]    io_outputs_0_combStage_translated_payload_size;
  wire                io_outputs_0_combStage_translated_payload_hasEarlyException;
  wire       [7:0]    io_outputs_0_combStage_translated_payload_earlyExceptionCode;
  wire       [1:0]    _zz_io_outputs_1_combStage_translated_payload_accessSize;
  wire                io_outputs_1_combStage_translated_valid;
  wire                io_outputs_1_combStage_translated_ready;
  wire       [31:0]   io_outputs_1_combStage_translated_payload_addr;
  wire       [31:0]   io_outputs_1_combStage_translated_payload_data;
  wire       [3:0]    io_outputs_1_combStage_translated_payload_be;
  wire       [3:0]    io_outputs_1_combStage_translated_payload_robPtr;
  wire       [1:0]    io_outputs_1_combStage_translated_payload_accessSize;
  wire                io_outputs_1_combStage_translated_payload_isFlush;
  wire                io_outputs_1_combStage_translated_payload_isIO;
  wire                io_outputs_1_combStage_translated_payload_hasEarlyException;
  wire       [7:0]    io_outputs_1_combStage_translated_payload_earlyExceptionCode;
  wire                LsuEU_LsuEuPlugin_hw_lqPushPort_fire;
  wire                StoreBufferPlugin_hw_pushPortInst_fire;
  wire                when_LsuEuPlugin_l141;
  wire                when_EuBasePlugin_l230_3;
  wire                LsuEU_LsuEuPlugin_logicPhase_executionCompletes;
  wire                LsuEU_LsuEuPlugin_logicPhase_completesSuccessfully;
  wire       [4:0]    _zz_when_Debug_l71_11;
  wire                when_Debug_l71_10;
  wire                when_EuBasePlugin_l300_3;
  reg                 s2_RobAlloc_ready_output;
  reg                 s1_Rename_ready_output;
  wire                when_Connection_l66_11;
  reg                 s0_Decode_ready_output;
  wire                when_Pipeline_l282;
  wire                when_Pipeline_l282_1;
  wire                when_Connection_l74;
  wire                when_Connection_l74_1;
  wire                when_Connection_l74_2;
  wire                _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid;
  reg        [2:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr;
  reg        [5:0]    _zz_when_AddressGenerationUnit_l215;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate;
  reg        [1:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc;
  reg        [5:0]    _zz_when_AddressGenerationUnit_l220;
  reg        [3:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad;
  reg                 _zz_when_AddressGenerationUnit_l220_1;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO;
  reg        [5:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_1;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_2;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_1;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_2;
  wire                when_AddressGenerationUnit_l215;
  wire                when_AddressGenerationUnit_l220;
  wire       [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_3;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_3;
  wire       [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_4;
  reg        [2:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_1;
  wire       [1:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask;
  reg        [3:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_1;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_input_ready;
  wire       [1:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize;
  wire                _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid_1;
  wire       [1:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid_2;
  reg        [2:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr_1;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_5;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_2;
  reg        [1:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2;
  reg        [3:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_2;
  reg        [5:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_basePhysReg;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate_1;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc_1;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc_1;
  reg        [3:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr_1;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad_1;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isStore;
  reg        [5:0]    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst_1;
  reg        [31:0]   _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_4;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush_1;
  reg                 _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO_1;
  wire                when_Stream_l477_5;
  wire                LoadQueuePlugin_logic_pushCmd_valid;
  wire                LoadQueuePlugin_logic_pushCmd_ready;
  wire       [3:0]    LoadQueuePlugin_logic_pushCmd_payload_robPtr;
  wire       [5:0]    LoadQueuePlugin_logic_pushCmd_payload_pdest;
  wire       [31:0]   LoadQueuePlugin_logic_pushCmd_payload_address;
  wire                LoadQueuePlugin_logic_pushCmd_payload_isIO;
  wire       [1:0]    LoadQueuePlugin_logic_pushCmd_payload_size;
  wire                LoadQueuePlugin_logic_pushCmd_payload_hasEarlyException;
  wire       [7:0]    LoadQueuePlugin_logic_pushCmd_payload_earlyExceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_0_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slots_0_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slots_0_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slots_0_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slots_0_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_0_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_0_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slots_0_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_0_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_1_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slots_1_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slots_1_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slots_1_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slots_1_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_1_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_1_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slots_1_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_1_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_1_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_1_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_1_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_2_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slots_2_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slots_2_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slots_2_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slots_2_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_2_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_2_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slots_2_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_2_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_2_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_2_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_2_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_3_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slots_3_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slots_3_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slots_3_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slots_3_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_3_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_3_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slots_3_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_3_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_3_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_3_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slots_3_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfo_valid;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfo_fromFwd;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfo_fromDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfo_fromMMIO;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfo_fromEarlyExc;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_completionInfo_data;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfo_hasFault;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_completionInfo_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromFwd;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromMMIO;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromEarlyExc;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_completionInfoReg_data;
  reg                 LoadQueuePlugin_logic_loadQueue_completionInfoReg_hasFault;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_completionInfoReg_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_0_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slotsNext_0_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_0_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_0_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_0_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_0_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_0_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_0_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_0_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_0_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_1_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slotsNext_1_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_1_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_1_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_1_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_1_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_1_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_1_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_1_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_1_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_2_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slotsNext_2_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_2_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_2_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_2_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_2_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_2_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_2_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_2_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_2_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_3_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_slotsNext_3_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_3_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_3_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_3_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_3_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_3_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_slotsNext_3_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_3_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_3_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_hit;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_data;
  reg                 LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_olderStoreHasUnknownAddress;
  reg                 LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_olderStoreDataNotReady;
  reg                 LoadQueuePlugin_logic_loadQueue_sbQueryRspValid;
  wire                LoadQueuePlugin_logic_loadQueue_flushInProgress;
  reg                 LoadQueuePlugin_logic_loadQueue_registeredFlush_valid;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr;
  wire                when_LoadQueuePlugin_l291;
  wire                LoadQueuePlugin_logic_loadQueue_canPush;
  wire       [3:0]    LoadQueuePlugin_logic_loadQueue_availableSlotsMask;
  wire       [3:0]    LoadQueuePlugin_logic_loadQueue_pushOh;
  wire                _zz_LoadQueuePlugin_logic_loadQueue_pushIdx;
  wire                _zz_LoadQueuePlugin_logic_loadQueue_pushIdx_1;
  wire                _zz_LoadQueuePlugin_logic_loadQueue_pushIdx_2;
  wire       [1:0]    LoadQueuePlugin_logic_loadQueue_pushIdx;
  wire                LoadQueuePlugin_logic_pushCmd_fire;
  wire       [3:0]    _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible;
  wire       [2:0]    _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_1;
  wire                _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_2;
  wire       [2:0]    _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_3;
  wire                LoadQueuePlugin_logic_loadQueue_headIsVisible;
  wire                LoadQueuePlugin_logic_loadQueue_headIsReadyForFwdQuery;
  wire                when_LoadQueuePlugin_l329;
  wire                when_LoadQueuePlugin_l335;
  wire                when_LoadQueuePlugin_l350;
  wire                LoadQueuePlugin_logic_loadQueue_headIsReadyToExecute;
  wire                LoadQueuePlugin_logic_loadQueue_shouldNotSendToMemory;
  reg        [1:0]    _zz_LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size;
  wire                LoadQueuePlugin_hw_dCacheLoadPort_cmd_fire;
  wire                LoadQueuePlugin_logic_loadQueue_mmioCmdFired;
  wire                LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead;
  wire                when_LoadQueuePlugin_l409;
  wire                LoadQueuePlugin_logic_loadQueue_popOnFwdHit;
  wire                LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess;
  wire                LoadQueuePlugin_logic_loadQueue_popOnEarlyException;
  wire                LoadQueuePlugin_logic_loadQueue_popRequest;
  reg                 LoadQueuePlugin_logic_loadQueue_completingHead_valid;
  reg        [31:0]   LoadQueuePlugin_logic_loadQueue_completingHead_address;
  reg        [1:0]    LoadQueuePlugin_logic_loadQueue_completingHead_size;
  reg        [3:0]    LoadQueuePlugin_logic_loadQueue_completingHead_robPtr;
  reg        [5:0]    LoadQueuePlugin_logic_loadQueue_completingHead_pdest;
  reg                 LoadQueuePlugin_logic_loadQueue_completingHead_isIO;
  reg                 LoadQueuePlugin_logic_loadQueue_completingHead_hasException;
  reg        [7:0]    LoadQueuePlugin_logic_loadQueue_completingHead_exceptionCode;
  reg                 LoadQueuePlugin_logic_loadQueue_completingHead_isWaitingForFwdRsp;
  reg                 LoadQueuePlugin_logic_loadQueue_completingHead_isStalledByDependency;
  reg                 LoadQueuePlugin_logic_loadQueue_completingHead_isReadyForDCache;
  reg                 LoadQueuePlugin_logic_loadQueue_completingHead_isWaitingForRsp;
  wire                when_LoadQueuePlugin_l478;
  wire                _zz_when_LoadQueuePlugin_l508;
  wire       [2:0]    _zz_when_LoadQueuePlugin_l508_1;
  wire                _zz_when_LoadQueuePlugin_l508_2;
  wire       [2:0]    _zz_when_LoadQueuePlugin_l508_3;
  wire                when_LoadQueuePlugin_l508;
  wire                _zz_when_LoadQueuePlugin_l508_4;
  wire       [2:0]    _zz_when_LoadQueuePlugin_l508_5;
  wire                _zz_when_LoadQueuePlugin_l508_6;
  wire       [2:0]    _zz_when_LoadQueuePlugin_l508_7;
  wire                when_LoadQueuePlugin_l508_1;
  wire                _zz_when_LoadQueuePlugin_l508_8;
  wire       [2:0]    _zz_when_LoadQueuePlugin_l508_9;
  wire                _zz_when_LoadQueuePlugin_l508_10;
  wire       [2:0]    _zz_when_LoadQueuePlugin_l508_11;
  wire                when_LoadQueuePlugin_l508_2;
  wire                _zz_when_LoadQueuePlugin_l508_12;
  wire       [2:0]    _zz_when_LoadQueuePlugin_l508_13;
  wire                _zz_when_LoadQueuePlugin_l508_14;
  wire       [2:0]    _zz_when_LoadQueuePlugin_l508_15;
  wire                when_LoadQueuePlugin_l508_3;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_0;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_1;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_2;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_3;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_4;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_5;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_6;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_7;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_8;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_9;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_10;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_11;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_12;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_13;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_14;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_15;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_16;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_17;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_18;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_19;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_20;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_21;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_22;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_23;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_24;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_25;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_26;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_27;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_28;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_29;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_30;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_31;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_32;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_33;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_34;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_35;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_36;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_37;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_38;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_39;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_40;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_41;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_42;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_43;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_44;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_45;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_46;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_47;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_48;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_49;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_50;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_51;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_52;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_53;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_54;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_55;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_56;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_57;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_58;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_59;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_60;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_61;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_62;
  reg        [31:0]   PhysicalRegFilePlugin_logic_regFile_63;
  wire                when_PhysicalRegFile_l130;
  wire       [63:0]   _zz_58;
  wire                when_PhysicalRegFile_l130_1;
  wire       [63:0]   _zz_59;
  wire                when_PhysicalRegFile_l130_2;
  wire       [63:0]   _zz_60;
  wire                when_PhysicalRegFile_l130_3;
  wire       [63:0]   _zz_61;
  wire                when_PhysicalRegFile_l130_4;
  wire       [63:0]   _zz_62;
  reg                 StoreBufferPlugin_logic_slots_0_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slots_0_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slots_0_data;
  reg        [3:0]    StoreBufferPlugin_logic_slots_0_be;
  reg        [3:0]    StoreBufferPlugin_logic_slots_0_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slots_0_accessSize;
  reg                 StoreBufferPlugin_logic_slots_0_isIO;
  reg                 StoreBufferPlugin_logic_slots_0_valid;
  reg                 StoreBufferPlugin_logic_slots_0_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slots_0_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slots_0_isCommitted;
  reg                 StoreBufferPlugin_logic_slots_0_sentCmd;
  reg                 StoreBufferPlugin_logic_slots_0_waitRsp;
  reg                 StoreBufferPlugin_logic_slots_0_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slots_0_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slots_0_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slots_1_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slots_1_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slots_1_data;
  reg        [3:0]    StoreBufferPlugin_logic_slots_1_be;
  reg        [3:0]    StoreBufferPlugin_logic_slots_1_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slots_1_accessSize;
  reg                 StoreBufferPlugin_logic_slots_1_isIO;
  reg                 StoreBufferPlugin_logic_slots_1_valid;
  reg                 StoreBufferPlugin_logic_slots_1_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slots_1_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slots_1_isCommitted;
  reg                 StoreBufferPlugin_logic_slots_1_sentCmd;
  reg                 StoreBufferPlugin_logic_slots_1_waitRsp;
  reg                 StoreBufferPlugin_logic_slots_1_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slots_1_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slots_1_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slots_2_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slots_2_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slots_2_data;
  reg        [3:0]    StoreBufferPlugin_logic_slots_2_be;
  reg        [3:0]    StoreBufferPlugin_logic_slots_2_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slots_2_accessSize;
  reg                 StoreBufferPlugin_logic_slots_2_isIO;
  reg                 StoreBufferPlugin_logic_slots_2_valid;
  reg                 StoreBufferPlugin_logic_slots_2_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slots_2_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slots_2_isCommitted;
  reg                 StoreBufferPlugin_logic_slots_2_sentCmd;
  reg                 StoreBufferPlugin_logic_slots_2_waitRsp;
  reg                 StoreBufferPlugin_logic_slots_2_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slots_2_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slots_2_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slots_3_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slots_3_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slots_3_data;
  reg        [3:0]    StoreBufferPlugin_logic_slots_3_be;
  reg        [3:0]    StoreBufferPlugin_logic_slots_3_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slots_3_accessSize;
  reg                 StoreBufferPlugin_logic_slots_3_isIO;
  reg                 StoreBufferPlugin_logic_slots_3_valid;
  reg                 StoreBufferPlugin_logic_slots_3_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slots_3_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slots_3_isCommitted;
  reg                 StoreBufferPlugin_logic_slots_3_sentCmd;
  reg                 StoreBufferPlugin_logic_slots_3_waitRsp;
  reg                 StoreBufferPlugin_logic_slots_3_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slots_3_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slots_3_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slotsAfterUpdates_0_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slotsAfterUpdates_0_data;
  reg        [3:0]    StoreBufferPlugin_logic_slotsAfterUpdates_0_be;
  reg        [3:0]    StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_valid;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_isCommitted;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slotsAfterUpdates_0_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slotsAfterUpdates_1_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slotsAfterUpdates_1_data;
  reg        [3:0]    StoreBufferPlugin_logic_slotsAfterUpdates_1_be;
  reg        [3:0]    StoreBufferPlugin_logic_slotsAfterUpdates_1_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_isIO;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_valid;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slotsAfterUpdates_1_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_isCommitted;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_sentCmd;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_waitRsp;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slotsAfterUpdates_1_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slotsAfterUpdates_2_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slotsAfterUpdates_2_data;
  reg        [3:0]    StoreBufferPlugin_logic_slotsAfterUpdates_2_be;
  reg        [3:0]    StoreBufferPlugin_logic_slotsAfterUpdates_2_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_isIO;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_valid;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slotsAfterUpdates_2_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_isCommitted;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_sentCmd;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_waitRsp;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slotsAfterUpdates_2_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slotsAfterUpdates_3_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slotsAfterUpdates_3_data;
  reg        [3:0]    StoreBufferPlugin_logic_slotsAfterUpdates_3_be;
  reg        [3:0]    StoreBufferPlugin_logic_slotsAfterUpdates_3_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_isIO;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_valid;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slotsAfterUpdates_3_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_isCommitted;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_sentCmd;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_waitRsp;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slotsAfterUpdates_3_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slotsNext_0_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slotsNext_0_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slotsNext_0_data;
  reg        [3:0]    StoreBufferPlugin_logic_slotsNext_0_be;
  reg        [3:0]    StoreBufferPlugin_logic_slotsNext_0_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slotsNext_0_accessSize;
  reg                 StoreBufferPlugin_logic_slotsNext_0_isIO;
  reg                 StoreBufferPlugin_logic_slotsNext_0_valid;
  reg                 StoreBufferPlugin_logic_slotsNext_0_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slotsNext_0_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slotsNext_0_isCommitted;
  reg                 StoreBufferPlugin_logic_slotsNext_0_sentCmd;
  reg                 StoreBufferPlugin_logic_slotsNext_0_waitRsp;
  reg                 StoreBufferPlugin_logic_slotsNext_0_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slotsNext_0_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slotsNext_0_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slotsNext_1_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slotsNext_1_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slotsNext_1_data;
  reg        [3:0]    StoreBufferPlugin_logic_slotsNext_1_be;
  reg        [3:0]    StoreBufferPlugin_logic_slotsNext_1_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slotsNext_1_accessSize;
  reg                 StoreBufferPlugin_logic_slotsNext_1_isIO;
  reg                 StoreBufferPlugin_logic_slotsNext_1_valid;
  reg                 StoreBufferPlugin_logic_slotsNext_1_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slotsNext_1_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slotsNext_1_isCommitted;
  reg                 StoreBufferPlugin_logic_slotsNext_1_sentCmd;
  reg                 StoreBufferPlugin_logic_slotsNext_1_waitRsp;
  reg                 StoreBufferPlugin_logic_slotsNext_1_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slotsNext_1_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slotsNext_1_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slotsNext_2_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slotsNext_2_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slotsNext_2_data;
  reg        [3:0]    StoreBufferPlugin_logic_slotsNext_2_be;
  reg        [3:0]    StoreBufferPlugin_logic_slotsNext_2_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slotsNext_2_accessSize;
  reg                 StoreBufferPlugin_logic_slotsNext_2_isIO;
  reg                 StoreBufferPlugin_logic_slotsNext_2_valid;
  reg                 StoreBufferPlugin_logic_slotsNext_2_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slotsNext_2_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slotsNext_2_isCommitted;
  reg                 StoreBufferPlugin_logic_slotsNext_2_sentCmd;
  reg                 StoreBufferPlugin_logic_slotsNext_2_waitRsp;
  reg                 StoreBufferPlugin_logic_slotsNext_2_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slotsNext_2_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slotsNext_2_refillSlotToWatch;
  reg                 StoreBufferPlugin_logic_slotsNext_3_isFlush;
  reg        [31:0]   StoreBufferPlugin_logic_slotsNext_3_addr;
  reg        [31:0]   StoreBufferPlugin_logic_slotsNext_3_data;
  reg        [3:0]    StoreBufferPlugin_logic_slotsNext_3_be;
  reg        [3:0]    StoreBufferPlugin_logic_slotsNext_3_robPtr;
  reg        [1:0]    StoreBufferPlugin_logic_slotsNext_3_accessSize;
  reg                 StoreBufferPlugin_logic_slotsNext_3_isIO;
  reg                 StoreBufferPlugin_logic_slotsNext_3_valid;
  reg                 StoreBufferPlugin_logic_slotsNext_3_hasEarlyException;
  reg        [7:0]    StoreBufferPlugin_logic_slotsNext_3_earlyExceptionCode;
  reg                 StoreBufferPlugin_logic_slotsNext_3_isCommitted;
  reg                 StoreBufferPlugin_logic_slotsNext_3_sentCmd;
  reg                 StoreBufferPlugin_logic_slotsNext_3_waitRsp;
  reg                 StoreBufferPlugin_logic_slotsNext_3_isWaitingForRefill;
  reg                 StoreBufferPlugin_logic_slotsNext_3_isWaitingForWb;
  reg        [7:0]    StoreBufferPlugin_logic_slotsNext_3_refillSlotToWatch;
  wire                StoreBufferPlugin_logic_flushInProgress;
  reg                 StoreBufferPlugin_logic_registeredFlush_valid;
  reg        [3:0]    StoreBufferPlugin_logic_registeredFlush_targetRobPtr;
  wire                StoreBufferPlugin_logic_validFall_0;
  wire                StoreBufferPlugin_logic_validFall_1;
  wire                StoreBufferPlugin_logic_validFall_2;
  wire                StoreBufferPlugin_logic_validFall_3;
  wire                StoreBufferPlugin_logic_canPush;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush;
  wire       [31:0]   _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_addr;
  wire       [31:0]   _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_data;
  wire       [3:0]    _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_be;
  wire       [3:0]    _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr;
  wire       [1:0]    _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize;
  wire                _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO;
  wire                _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException;
  wire       [7:0]    _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode;
  wire       [3:0]    _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                StoreBufferPlugin_logic_sharedWriteCond;
  wire                StoreBufferPlugin_logic_canPopNormalOp;
  wire                StoreBufferPlugin_logic_canPopFlushOp;
  wire                StoreBufferPlugin_logic_canPopMMIOOp;
  wire                when_StoreBufferPlugin_l316;
  wire                StoreBufferPlugin_logic_canSendToDCache;
  wire                StoreBufferPlugin_logic_dcacheCmdFired;
  wire                StoreBufferPlugin_logic_mmioCmdFired;
  wire                StoreBufferPlugin_logic_dcacheResponseForHead;
  wire                StoreBufferPlugin_logic_mmioResponseForHead;
  wire       [5:0]    _zz_when_Debug_l71_12;
  wire                when_Debug_l71_11;
  wire                StoreBufferPlugin_logic_waitedRefillIsDone;
  wire                when_StoreBufferPlugin_l474;
  reg        [3:0]    StoreBufferPlugin_logic_commitUpdateInfo_validMask;
  reg                 _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask;
  wire                when_StoreBufferPlugin_l498;
  wire                when_StoreBufferPlugin_l504;
  reg                 _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_1;
  wire                when_StoreBufferPlugin_l498_1;
  wire                when_StoreBufferPlugin_l504_1;
  reg                 _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_2;
  wire                when_StoreBufferPlugin_l498_2;
  wire                when_StoreBufferPlugin_l504_2;
  reg                 _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_3;
  wire                when_StoreBufferPlugin_l498_3;
  wire                when_StoreBufferPlugin_l504_3;
  reg        [3:0]    StoreBufferPlugin_logic_registeredCommitUpdate_validMask;
  wire                _zz_when_StoreBufferPlugin_l525;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l525_1;
  wire                _zz_when_StoreBufferPlugin_l525_2;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l525_3;
  wire                when_StoreBufferPlugin_l525;
  wire                when_StoreBufferPlugin_l533;
  wire                when_StoreBufferPlugin_l529;
  wire                _zz_when_StoreBufferPlugin_l525_4;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l525_5;
  wire                _zz_when_StoreBufferPlugin_l525_6;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l525_7;
  wire                when_StoreBufferPlugin_l525_1;
  wire                when_StoreBufferPlugin_l533_1;
  wire                when_StoreBufferPlugin_l529_1;
  wire                _zz_when_StoreBufferPlugin_l525_8;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l525_9;
  wire                _zz_when_StoreBufferPlugin_l525_10;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l525_11;
  wire                when_StoreBufferPlugin_l525_2;
  wire                when_StoreBufferPlugin_l533_2;
  wire                when_StoreBufferPlugin_l529_2;
  wire                _zz_when_StoreBufferPlugin_l525_12;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l525_13;
  wire                _zz_when_StoreBufferPlugin_l525_14;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l525_15;
  wire                when_StoreBufferPlugin_l525_3;
  wire                when_StoreBufferPlugin_l533_3;
  wire                when_StoreBufferPlugin_l529_3;
  wire                when_StoreBufferPlugin_l540;
  wire                StoreBufferPlugin_logic_operationDone;
  reg                 StoreBufferPlugin_logic_popRequest;
  wire                when_StoreBufferPlugin_l555;
  wire                when_StoreBufferPlugin_l576;
  wire       [3:0]    StoreBufferPlugin_logic_forwardingLogic_loadMask;
  reg        [3:0]    _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask;
  wire       [1:0]    _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_1;
  wire       [31:0]   StoreBufferPlugin_logic_forwardingLogic_bypassInitial_data;
  wire       [3:0]    StoreBufferPlugin_logic_forwardingLogic_bypassInitial_hitMask;
  reg        [31:0]   _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data;
  reg        [3:0]    _zz_when_StoreBufferPlugin_l640;
  wire                _zz_when_StoreBufferPlugin_l631;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l631_1;
  wire                _zz_when_StoreBufferPlugin_l631_2;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l631_3;
  wire                when_StoreBufferPlugin_l631;
  wire                _zz_when_StoreBufferPlugin_l638;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l638_1;
  wire                _zz_when_StoreBufferPlugin_l638_2;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l638_3;
  wire                when_StoreBufferPlugin_l638;
  wire                when_StoreBufferPlugin_l640;
  wire                when_StoreBufferPlugin_l640_1;
  wire                when_StoreBufferPlugin_l640_2;
  wire                when_StoreBufferPlugin_l640_3;
  reg        [31:0]   _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_1;
  reg        [3:0]    _zz_when_StoreBufferPlugin_l640_1;
  wire                _zz_when_StoreBufferPlugin_l631_4;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l631_5;
  wire                _zz_when_StoreBufferPlugin_l631_6;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l631_7;
  wire                when_StoreBufferPlugin_l631_1;
  wire                _zz_when_StoreBufferPlugin_l638_4;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l638_5;
  wire                _zz_when_StoreBufferPlugin_l638_6;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l638_7;
  wire                when_StoreBufferPlugin_l638_1;
  wire                when_StoreBufferPlugin_l640_4;
  wire                when_StoreBufferPlugin_l640_5;
  wire                when_StoreBufferPlugin_l640_6;
  wire                when_StoreBufferPlugin_l640_7;
  reg        [31:0]   _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_2;
  reg        [3:0]    _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask;
  wire                _zz_when_StoreBufferPlugin_l631_8;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l631_9;
  wire                _zz_when_StoreBufferPlugin_l631_10;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l631_11;
  wire                when_StoreBufferPlugin_l631_2;
  wire                _zz_when_StoreBufferPlugin_l638_8;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l638_9;
  wire                _zz_when_StoreBufferPlugin_l638_10;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l638_11;
  wire                when_StoreBufferPlugin_l638_2;
  wire                when_StoreBufferPlugin_l640_8;
  wire                when_StoreBufferPlugin_l640_9;
  wire                when_StoreBufferPlugin_l640_10;
  wire                when_StoreBufferPlugin_l640_11;
  reg        [31:0]   StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data;
  reg        [3:0]    StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask;
  wire                _zz_when_StoreBufferPlugin_l631_12;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l631_13;
  wire                _zz_when_StoreBufferPlugin_l631_14;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l631_15;
  wire                when_StoreBufferPlugin_l631_3;
  wire                _zz_when_StoreBufferPlugin_l638_12;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l638_13;
  wire                _zz_when_StoreBufferPlugin_l638_14;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l638_15;
  wire                when_StoreBufferPlugin_l638_3;
  wire                when_StoreBufferPlugin_l640_12;
  wire                when_StoreBufferPlugin_l640_13;
  wire                when_StoreBufferPlugin_l640_14;
  wire                when_StoreBufferPlugin_l640_15;
  wire                StoreBufferPlugin_logic_forwardingLogic_allRequiredBytesHit;
  reg                 StoreBufferPlugin_logic_forwardingLogic_dataNotReadyStall;
  reg                 StoreBufferPlugin_logic_forwardingLogic_hasOlderOverlappingStore;
  wire                when_StoreBufferPlugin_l672;
  wire                _zz_when_StoreBufferPlugin_l678;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l678_1;
  wire                _zz_when_StoreBufferPlugin_l678_2;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l678_3;
  wire       [29:0]   _zz_when_StoreBufferPlugin_l678_4;
  wire       [29:0]   _zz_when_StoreBufferPlugin_l678_5;
  wire                when_StoreBufferPlugin_l678;
  wire                when_StoreBufferPlugin_l681;
  wire                when_StoreBufferPlugin_l672_1;
  wire                _zz_when_StoreBufferPlugin_l678_6;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l678_7;
  wire                _zz_when_StoreBufferPlugin_l678_8;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l678_9;
  wire       [29:0]   _zz_when_StoreBufferPlugin_l678_10;
  wire       [29:0]   _zz_when_StoreBufferPlugin_l678_11;
  wire                when_StoreBufferPlugin_l678_1;
  wire                when_StoreBufferPlugin_l681_1;
  wire                when_StoreBufferPlugin_l672_2;
  wire                _zz_when_StoreBufferPlugin_l678_12;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l678_13;
  wire                _zz_when_StoreBufferPlugin_l678_14;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l678_15;
  wire       [29:0]   _zz_when_StoreBufferPlugin_l678_16;
  wire       [29:0]   _zz_when_StoreBufferPlugin_l678_17;
  wire                when_StoreBufferPlugin_l678_2;
  wire                when_StoreBufferPlugin_l681_2;
  wire                when_StoreBufferPlugin_l672_3;
  wire                _zz_when_StoreBufferPlugin_l678_18;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l678_19;
  wire                _zz_when_StoreBufferPlugin_l678_20;
  wire       [2:0]    _zz_when_StoreBufferPlugin_l678_21;
  wire       [29:0]   _zz_when_StoreBufferPlugin_l678_22;
  wire       [29:0]   _zz_when_StoreBufferPlugin_l678_23;
  wire                when_StoreBufferPlugin_l678_3;
  wire                when_StoreBufferPlugin_l681_3;
  wire                StoreBufferPlugin_logic_forwardingLogic_insufficientCoverageStall;
  wire                StoreBufferPlugin_logic_bypassResult_hit;
  wire       [31:0]   StoreBufferPlugin_logic_bypassResult_data;
  wire       [3:0]    StoreBufferPlugin_logic_bypassResult_hitMask;
  reg        [3:0]    _zz_StoreBufferPlugin_logic_loadQueryBe;
  wire       [1:0]    _zz_StoreBufferPlugin_logic_loadQueryBe_1;
  wire       [3:0]    StoreBufferPlugin_logic_loadQueryBe;
  wire       [31:0]   StoreBufferPlugin_logic_bypassInitial_data;
  wire       [3:0]    StoreBufferPlugin_logic_bypassInitial_hitMask;
  reg        [31:0]   _zz_StoreBufferPlugin_logic_finalBypassResult_data;
  reg        [3:0]    _zz_when_StoreBufferPlugin_l742;
  wire                when_StoreBufferPlugin_l735;
  wire                when_StoreBufferPlugin_l740;
  wire                when_StoreBufferPlugin_l742;
  wire                when_StoreBufferPlugin_l742_1;
  wire                when_StoreBufferPlugin_l742_2;
  wire                when_StoreBufferPlugin_l742_3;
  reg        [31:0]   _zz_StoreBufferPlugin_logic_finalBypassResult_data_1;
  reg        [3:0]    _zz_when_StoreBufferPlugin_l742_1;
  wire                when_StoreBufferPlugin_l735_1;
  wire                when_StoreBufferPlugin_l740_1;
  wire                when_StoreBufferPlugin_l742_4;
  wire                when_StoreBufferPlugin_l742_5;
  wire                when_StoreBufferPlugin_l742_6;
  wire                when_StoreBufferPlugin_l742_7;
  reg        [31:0]   _zz_StoreBufferPlugin_logic_finalBypassResult_data_2;
  reg        [3:0]    _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask;
  wire                when_StoreBufferPlugin_l735_2;
  wire                when_StoreBufferPlugin_l740_2;
  wire                when_StoreBufferPlugin_l742_8;
  wire                when_StoreBufferPlugin_l742_9;
  wire                when_StoreBufferPlugin_l742_10;
  wire                when_StoreBufferPlugin_l742_11;
  reg        [31:0]   StoreBufferPlugin_logic_finalBypassResult_data;
  reg        [3:0]    StoreBufferPlugin_logic_finalBypassResult_hitMask;
  wire                when_StoreBufferPlugin_l735_3;
  wire                when_StoreBufferPlugin_l740_3;
  wire                when_StoreBufferPlugin_l742_12;
  wire                when_StoreBufferPlugin_l742_13;
  wire                when_StoreBufferPlugin_l742_14;
  wire                when_StoreBufferPlugin_l742_15;
  wire                StoreBufferPlugin_logic_overallBypassHit;
  wire       [63:0]   BusyTablePlugin_logic_busyTableNext;
  reg                 FetchPipelinePlugin_logic_retryIdCounter_willIncrement;
  wire                FetchPipelinePlugin_logic_retryIdCounter_willClear;
  reg        [1:0]    FetchPipelinePlugin_logic_retryIdCounter_valueNext;
  reg        [1:0]    FetchPipelinePlugin_logic_retryIdCounter_value;
  wire                FetchPipelinePlugin_logic_retryIdCounter_willOverflowIfInc;
  wire                FetchPipelinePlugin_logic_retryIdCounter_willOverflow;
  reg                 FetchPipelinePlugin_logic_doRetryFlush;
  wire                s1_PC_Gen_valid;
  reg                 _zz_s2_ICache_Access_valid;
  reg                 s2_ICache_Access_valid;
  reg                 _zz_s4_Predecode_valid;
  wire                s3_ICache_Wait_valid;
  reg                 s4_Predecode_valid;
  wire                FetchPipelinePlugin_logic_hardRedirect_valid;
  wire       [31:0]   FetchPipelinePlugin_logic_hardRedirect_payload;
  wire                FetchPipelinePlugin_logic_doAnyFlush;
  wire                io_pop_fire;
  reg                 FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_incrementIt;
  reg                 FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_decrementIt;
  wire       [2:0]    FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_valueNext;
  reg        [2:0]    FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value;
  wire                FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_mayOverflow;
  wire                FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_mayUnderflow;
  wire                FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willOverflowIfInc;
  wire                FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willOverflow;
  wire                FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willUnderflowIfDec;
  wire                FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willUnderflow;
  reg        [2:0]    FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_finalIncrement;
  wire                when_Utils_l767;
  wire                when_Utils_l769;
  reg                 FetchPipelinePlugin_logic_isDrainingCacheRspReg;
  wire                when_FetchPipelinePlugin2_l289;
  reg                 FetchPipelinePlugin_logic_retryCmd_lock;
  reg        [31:0]   FetchPipelinePlugin_logic_retryCmd_pc;
  reg        [1:0]    FetchPipelinePlugin_logic_retryCmd_id;
  reg        [31:0]   FetchPipelinePlugin_logic_s1_logic_fetchPcReg;
  reg        [1:0]    FetchPipelinePlugin_logic_s1_logic_lastRetryIdReg;
  wire                FetchPipelinePlugin_logic_s1_logic_needRedo;
  wire       [31:0]   FetchPipelinePlugin_logic_s1_logic_rawPcToUse;
  wire       [31:0]   FetchPipelinePlugin_logic_s1_logic_nextLinePc;
  wire       [31:0]   _zz_FetchPipelinePlugin_logic_s1_logic_fetchPcReg;
  wire                s1_PC_Gen_isFiring;
  wire                when_FetchPipelinePlugin2_l361;
  wire                when_FetchPipelinePlugin2_l367;
  wire                FetchPipelinePlugin_logic_s1_logic_fetchDisabled;
  wire                when_FetchPipelinePlugin2_l380;
  wire                s1_PC_Gen_haltRequest_FetchPipelinePlugin2_l381;
  wire                s2_ICache_Access_isFiring;
  wire       [31:0]   FetchPipelinePlugin_logic_s2_logic_cmdPayload_address;
  wire       [7:0]    FetchPipelinePlugin_logic_s2_logic_cmdPayload_transactionId;
  wire                s4_Predecode_isFiring;
  wire                FetchPipelinePlugin_logic_s4_logic_handleRsp;
  wire                FetchPipelinePlugin_logic_s4_logic_hasHigherPriorityStuff;
  wire                FetchPipelinePlugin_logic_s4_logic_backpressureRedo;
  wire                when_FetchPipelinePlugin2_l442;
  wire       [27:0]   _zz_70;
  wire                when_FetchPipelinePlugin2_l458;
  wire                when_FetchPipelinePlugin2_l467;
  wire                when_FetchPipelinePlugin2_l476;
  wire                when_FetchPipelinePlugin2_l481;
  wire                _zz_io_push_payload_predecodeInfos_0_isBranch;
  wire                _zz_io_push_payload_predecodeInfos_1_isBranch;
  wire                _zz_io_push_payload_predecodeInfos_2_isBranch;
  wire                _zz_io_push_payload_predecodeInfos_3_isBranch;
  wire       [2:0]    _zz_io_push_payload_numValidInstructions;
  wire       [1:0]    _zz_io_push_payload_startInstructionIndex;
  wire       [31:0]   _zz_io_push_payload_numValidInstructions_1;
  wire       [1:0]    _zz_io_push_payload_numValidInstructions_2;
  wire                s4_Predecode_haltRequest_FetchPipelinePlugin2_l505;
  wire                io_push_fire;
  wire                io_fetchGroupIn_fire;
  wire                _zz_71;
  wire                _zz_s2_ICache_Access_isFlushingRoot;
  wire                _zz_s3_ICache_Wait_isFlushingRoot;
  reg                 s2_ICache_Access_ready_output;
  wire                when_Connection_l66_12;
  reg                 s1_PC_Gen_ready_output;
  wire                when_Pipeline_l282_2;
  wire                when_Pipeline_l282_3;
  wire                when_Connection_l74_3;
  wire                when_Connection_l74_4;
  wire       [0:0]    DataCachePlugin_logic_load_hits;
  wire                DataCachePlugin_logic_load_hit;
  wire                DataCachePlugin_logic_load_hits_bools_0;
  wire       [0:0]    _zz_DataCachePlugin_logic_load_oh;
  wire       [0:0]    DataCachePlugin_logic_load_oh;
  wire       [0:0]    DataCachePlugin_logic_load_ohHistory_0;
  wire       [0:0]    DataCachePlugin_logic_load_ohHistory_1;
  wire       [0:0]    DataCachePlugin_logic_load_ohHistory_2;
  wire       [0:0]    _zz_DataCachePlugin_logic_load_ohHistory_0;
  reg        [0:0]    _zz_DataCachePlugin_logic_load_ohHistory_1;
  reg        [0:0]    _zz_DataCachePlugin_logic_load_ohHistory_2;
  reg        [1:0]    _zz_ROBPlugin_aggregatedFlushSignal_payload_reason;
  reg        [3:0]    _zz_ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr;
  reg                 ICachePlugin_axiMaster_ar_valid;
  wire                ICachePlugin_axiMaster_ar_ready;
  reg        [31:0]   ICachePlugin_axiMaster_ar_payload_addr;
  wire       [3:0]    ICachePlugin_axiMaster_ar_payload_id;
  reg        [7:0]    ICachePlugin_axiMaster_ar_payload_len;
  reg        [2:0]    ICachePlugin_axiMaster_ar_payload_size;
  reg        [1:0]    ICachePlugin_axiMaster_ar_payload_burst;
  wire                ICachePlugin_axiMaster_r_valid;
  reg                 ICachePlugin_axiMaster_r_ready;
  wire       [31:0]   ICachePlugin_axiMaster_r_payload_data;
  wire       [3:0]    ICachePlugin_axiMaster_r_payload_id;
  wire       [1:0]    ICachePlugin_axiMaster_r_payload_resp;
  wire                ICachePlugin_axiMaster_r_payload_last;
  wire                CoreMemSysPlugin_logic_roMasters_0_aw_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_aw_ready;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_aw_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_aw_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_aw_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_aw_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_aw_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_w_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_w_ready;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_w_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_w_payload_strb;
  wire                CoreMemSysPlugin_logic_roMasters_0_w_payload_last;
  wire                CoreMemSysPlugin_logic_roMasters_0_b_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_b_ready;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_b_payload_id;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_b_payload_resp;
  wire                CoreMemSysPlugin_logic_roMasters_0_ar_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_ar_ready;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_ar_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_ar_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_ar_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_ar_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_ar_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_r_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_r_ready;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_r_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_r_payload_id;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_r_payload_resp;
  wire                CoreMemSysPlugin_logic_roMasters_0_r_payload_last;
  wire                when_CheckpointManagerPlugin_l117;
  wire                when_CheckpointManagerPlugin_l121;
  reg                 ICachePlugin_logic_storage_valids_0_0;
  reg                 ICachePlugin_logic_storage_valids_0_1;
  reg                 ICachePlugin_logic_storage_valids_1_0;
  reg                 ICachePlugin_logic_storage_valids_1_1;
  reg                 ICachePlugin_logic_storage_valids_2_0;
  reg                 ICachePlugin_logic_storage_valids_2_1;
  reg                 ICachePlugin_logic_storage_valids_3_0;
  reg                 ICachePlugin_logic_storage_valids_3_1;
  reg                 ICachePlugin_logic_storage_valids_4_0;
  reg                 ICachePlugin_logic_storage_valids_4_1;
  reg                 ICachePlugin_logic_storage_valids_5_0;
  reg                 ICachePlugin_logic_storage_valids_5_1;
  reg                 ICachePlugin_logic_storage_valids_6_0;
  reg                 ICachePlugin_logic_storage_valids_6_1;
  reg                 ICachePlugin_logic_storage_valids_7_0;
  reg                 ICachePlugin_logic_storage_valids_7_1;
  reg                 ICachePlugin_logic_storage_valids_8_0;
  reg                 ICachePlugin_logic_storage_valids_8_1;
  reg                 ICachePlugin_logic_storage_valids_9_0;
  reg                 ICachePlugin_logic_storage_valids_9_1;
  reg                 ICachePlugin_logic_storage_valids_10_0;
  reg                 ICachePlugin_logic_storage_valids_10_1;
  reg                 ICachePlugin_logic_storage_valids_11_0;
  reg                 ICachePlugin_logic_storage_valids_11_1;
  reg                 ICachePlugin_logic_storage_valids_12_0;
  reg                 ICachePlugin_logic_storage_valids_12_1;
  reg                 ICachePlugin_logic_storage_valids_13_0;
  reg                 ICachePlugin_logic_storage_valids_13_1;
  reg                 ICachePlugin_logic_storage_valids_14_0;
  reg                 ICachePlugin_logic_storage_valids_14_1;
  reg                 ICachePlugin_logic_storage_valids_15_0;
  reg                 ICachePlugin_logic_storage_valids_15_1;
  reg                 ICachePlugin_logic_storage_valids_16_0;
  reg                 ICachePlugin_logic_storage_valids_16_1;
  reg                 ICachePlugin_logic_storage_valids_17_0;
  reg                 ICachePlugin_logic_storage_valids_17_1;
  reg                 ICachePlugin_logic_storage_valids_18_0;
  reg                 ICachePlugin_logic_storage_valids_18_1;
  reg                 ICachePlugin_logic_storage_valids_19_0;
  reg                 ICachePlugin_logic_storage_valids_19_1;
  reg                 ICachePlugin_logic_storage_valids_20_0;
  reg                 ICachePlugin_logic_storage_valids_20_1;
  reg                 ICachePlugin_logic_storage_valids_21_0;
  reg                 ICachePlugin_logic_storage_valids_21_1;
  reg                 ICachePlugin_logic_storage_valids_22_0;
  reg                 ICachePlugin_logic_storage_valids_22_1;
  reg                 ICachePlugin_logic_storage_valids_23_0;
  reg                 ICachePlugin_logic_storage_valids_23_1;
  reg                 ICachePlugin_logic_storage_valids_24_0;
  reg                 ICachePlugin_logic_storage_valids_24_1;
  reg                 ICachePlugin_logic_storage_valids_25_0;
  reg                 ICachePlugin_logic_storage_valids_25_1;
  reg                 ICachePlugin_logic_storage_valids_26_0;
  reg                 ICachePlugin_logic_storage_valids_26_1;
  reg                 ICachePlugin_logic_storage_valids_27_0;
  reg                 ICachePlugin_logic_storage_valids_27_1;
  reg                 ICachePlugin_logic_storage_valids_28_0;
  reg                 ICachePlugin_logic_storage_valids_28_1;
  reg                 ICachePlugin_logic_storage_valids_29_0;
  reg                 ICachePlugin_logic_storage_valids_29_1;
  reg                 ICachePlugin_logic_storage_valids_30_0;
  reg                 ICachePlugin_logic_storage_valids_30_1;
  reg                 ICachePlugin_logic_storage_valids_31_0;
  reg                 ICachePlugin_logic_storage_valids_31_1;
  reg                 ICachePlugin_logic_storage_valids_32_0;
  reg                 ICachePlugin_logic_storage_valids_32_1;
  reg                 ICachePlugin_logic_storage_valids_33_0;
  reg                 ICachePlugin_logic_storage_valids_33_1;
  reg                 ICachePlugin_logic_storage_valids_34_0;
  reg                 ICachePlugin_logic_storage_valids_34_1;
  reg                 ICachePlugin_logic_storage_valids_35_0;
  reg                 ICachePlugin_logic_storage_valids_35_1;
  reg                 ICachePlugin_logic_storage_valids_36_0;
  reg                 ICachePlugin_logic_storage_valids_36_1;
  reg                 ICachePlugin_logic_storage_valids_37_0;
  reg                 ICachePlugin_logic_storage_valids_37_1;
  reg                 ICachePlugin_logic_storage_valids_38_0;
  reg                 ICachePlugin_logic_storage_valids_38_1;
  reg                 ICachePlugin_logic_storage_valids_39_0;
  reg                 ICachePlugin_logic_storage_valids_39_1;
  reg                 ICachePlugin_logic_storage_valids_40_0;
  reg                 ICachePlugin_logic_storage_valids_40_1;
  reg                 ICachePlugin_logic_storage_valids_41_0;
  reg                 ICachePlugin_logic_storage_valids_41_1;
  reg                 ICachePlugin_logic_storage_valids_42_0;
  reg                 ICachePlugin_logic_storage_valids_42_1;
  reg                 ICachePlugin_logic_storage_valids_43_0;
  reg                 ICachePlugin_logic_storage_valids_43_1;
  reg                 ICachePlugin_logic_storage_valids_44_0;
  reg                 ICachePlugin_logic_storage_valids_44_1;
  reg                 ICachePlugin_logic_storage_valids_45_0;
  reg                 ICachePlugin_logic_storage_valids_45_1;
  reg                 ICachePlugin_logic_storage_valids_46_0;
  reg                 ICachePlugin_logic_storage_valids_46_1;
  reg                 ICachePlugin_logic_storage_valids_47_0;
  reg                 ICachePlugin_logic_storage_valids_47_1;
  reg                 ICachePlugin_logic_storage_valids_48_0;
  reg                 ICachePlugin_logic_storage_valids_48_1;
  reg                 ICachePlugin_logic_storage_valids_49_0;
  reg                 ICachePlugin_logic_storage_valids_49_1;
  reg                 ICachePlugin_logic_storage_valids_50_0;
  reg                 ICachePlugin_logic_storage_valids_50_1;
  reg                 ICachePlugin_logic_storage_valids_51_0;
  reg                 ICachePlugin_logic_storage_valids_51_1;
  reg                 ICachePlugin_logic_storage_valids_52_0;
  reg                 ICachePlugin_logic_storage_valids_52_1;
  reg                 ICachePlugin_logic_storage_valids_53_0;
  reg                 ICachePlugin_logic_storage_valids_53_1;
  reg                 ICachePlugin_logic_storage_valids_54_0;
  reg                 ICachePlugin_logic_storage_valids_54_1;
  reg                 ICachePlugin_logic_storage_valids_55_0;
  reg                 ICachePlugin_logic_storage_valids_55_1;
  reg                 ICachePlugin_logic_storage_valids_56_0;
  reg                 ICachePlugin_logic_storage_valids_56_1;
  reg                 ICachePlugin_logic_storage_valids_57_0;
  reg                 ICachePlugin_logic_storage_valids_57_1;
  reg                 ICachePlugin_logic_storage_valids_58_0;
  reg                 ICachePlugin_logic_storage_valids_58_1;
  reg                 ICachePlugin_logic_storage_valids_59_0;
  reg                 ICachePlugin_logic_storage_valids_59_1;
  reg                 ICachePlugin_logic_storage_valids_60_0;
  reg                 ICachePlugin_logic_storage_valids_60_1;
  reg                 ICachePlugin_logic_storage_valids_61_0;
  reg                 ICachePlugin_logic_storage_valids_61_1;
  reg                 ICachePlugin_logic_storage_valids_62_0;
  reg                 ICachePlugin_logic_storage_valids_62_1;
  reg                 ICachePlugin_logic_storage_valids_63_0;
  reg                 ICachePlugin_logic_storage_valids_63_1;
  reg                 ICachePlugin_logic_storage_valids_64_0;
  reg                 ICachePlugin_logic_storage_valids_64_1;
  reg                 ICachePlugin_logic_storage_valids_65_0;
  reg                 ICachePlugin_logic_storage_valids_65_1;
  reg                 ICachePlugin_logic_storage_valids_66_0;
  reg                 ICachePlugin_logic_storage_valids_66_1;
  reg                 ICachePlugin_logic_storage_valids_67_0;
  reg                 ICachePlugin_logic_storage_valids_67_1;
  reg                 ICachePlugin_logic_storage_valids_68_0;
  reg                 ICachePlugin_logic_storage_valids_68_1;
  reg                 ICachePlugin_logic_storage_valids_69_0;
  reg                 ICachePlugin_logic_storage_valids_69_1;
  reg                 ICachePlugin_logic_storage_valids_70_0;
  reg                 ICachePlugin_logic_storage_valids_70_1;
  reg                 ICachePlugin_logic_storage_valids_71_0;
  reg                 ICachePlugin_logic_storage_valids_71_1;
  reg                 ICachePlugin_logic_storage_valids_72_0;
  reg                 ICachePlugin_logic_storage_valids_72_1;
  reg                 ICachePlugin_logic_storage_valids_73_0;
  reg                 ICachePlugin_logic_storage_valids_73_1;
  reg                 ICachePlugin_logic_storage_valids_74_0;
  reg                 ICachePlugin_logic_storage_valids_74_1;
  reg                 ICachePlugin_logic_storage_valids_75_0;
  reg                 ICachePlugin_logic_storage_valids_75_1;
  reg                 ICachePlugin_logic_storage_valids_76_0;
  reg                 ICachePlugin_logic_storage_valids_76_1;
  reg                 ICachePlugin_logic_storage_valids_77_0;
  reg                 ICachePlugin_logic_storage_valids_77_1;
  reg                 ICachePlugin_logic_storage_valids_78_0;
  reg                 ICachePlugin_logic_storage_valids_78_1;
  reg                 ICachePlugin_logic_storage_valids_79_0;
  reg                 ICachePlugin_logic_storage_valids_79_1;
  reg                 ICachePlugin_logic_storage_valids_80_0;
  reg                 ICachePlugin_logic_storage_valids_80_1;
  reg                 ICachePlugin_logic_storage_valids_81_0;
  reg                 ICachePlugin_logic_storage_valids_81_1;
  reg                 ICachePlugin_logic_storage_valids_82_0;
  reg                 ICachePlugin_logic_storage_valids_82_1;
  reg                 ICachePlugin_logic_storage_valids_83_0;
  reg                 ICachePlugin_logic_storage_valids_83_1;
  reg                 ICachePlugin_logic_storage_valids_84_0;
  reg                 ICachePlugin_logic_storage_valids_84_1;
  reg                 ICachePlugin_logic_storage_valids_85_0;
  reg                 ICachePlugin_logic_storage_valids_85_1;
  reg                 ICachePlugin_logic_storage_valids_86_0;
  reg                 ICachePlugin_logic_storage_valids_86_1;
  reg                 ICachePlugin_logic_storage_valids_87_0;
  reg                 ICachePlugin_logic_storage_valids_87_1;
  reg                 ICachePlugin_logic_storage_valids_88_0;
  reg                 ICachePlugin_logic_storage_valids_88_1;
  reg                 ICachePlugin_logic_storage_valids_89_0;
  reg                 ICachePlugin_logic_storage_valids_89_1;
  reg                 ICachePlugin_logic_storage_valids_90_0;
  reg                 ICachePlugin_logic_storage_valids_90_1;
  reg                 ICachePlugin_logic_storage_valids_91_0;
  reg                 ICachePlugin_logic_storage_valids_91_1;
  reg                 ICachePlugin_logic_storage_valids_92_0;
  reg                 ICachePlugin_logic_storage_valids_92_1;
  reg                 ICachePlugin_logic_storage_valids_93_0;
  reg                 ICachePlugin_logic_storage_valids_93_1;
  reg                 ICachePlugin_logic_storage_valids_94_0;
  reg                 ICachePlugin_logic_storage_valids_94_1;
  reg                 ICachePlugin_logic_storage_valids_95_0;
  reg                 ICachePlugin_logic_storage_valids_95_1;
  reg                 ICachePlugin_logic_storage_valids_96_0;
  reg                 ICachePlugin_logic_storage_valids_96_1;
  reg                 ICachePlugin_logic_storage_valids_97_0;
  reg                 ICachePlugin_logic_storage_valids_97_1;
  reg                 ICachePlugin_logic_storage_valids_98_0;
  reg                 ICachePlugin_logic_storage_valids_98_1;
  reg                 ICachePlugin_logic_storage_valids_99_0;
  reg                 ICachePlugin_logic_storage_valids_99_1;
  reg                 ICachePlugin_logic_storage_valids_100_0;
  reg                 ICachePlugin_logic_storage_valids_100_1;
  reg                 ICachePlugin_logic_storage_valids_101_0;
  reg                 ICachePlugin_logic_storage_valids_101_1;
  reg                 ICachePlugin_logic_storage_valids_102_0;
  reg                 ICachePlugin_logic_storage_valids_102_1;
  reg                 ICachePlugin_logic_storage_valids_103_0;
  reg                 ICachePlugin_logic_storage_valids_103_1;
  reg                 ICachePlugin_logic_storage_valids_104_0;
  reg                 ICachePlugin_logic_storage_valids_104_1;
  reg                 ICachePlugin_logic_storage_valids_105_0;
  reg                 ICachePlugin_logic_storage_valids_105_1;
  reg                 ICachePlugin_logic_storage_valids_106_0;
  reg                 ICachePlugin_logic_storage_valids_106_1;
  reg                 ICachePlugin_logic_storage_valids_107_0;
  reg                 ICachePlugin_logic_storage_valids_107_1;
  reg                 ICachePlugin_logic_storage_valids_108_0;
  reg                 ICachePlugin_logic_storage_valids_108_1;
  reg                 ICachePlugin_logic_storage_valids_109_0;
  reg                 ICachePlugin_logic_storage_valids_109_1;
  reg                 ICachePlugin_logic_storage_valids_110_0;
  reg                 ICachePlugin_logic_storage_valids_110_1;
  reg                 ICachePlugin_logic_storage_valids_111_0;
  reg                 ICachePlugin_logic_storage_valids_111_1;
  reg                 ICachePlugin_logic_storage_valids_112_0;
  reg                 ICachePlugin_logic_storage_valids_112_1;
  reg                 ICachePlugin_logic_storage_valids_113_0;
  reg                 ICachePlugin_logic_storage_valids_113_1;
  reg                 ICachePlugin_logic_storage_valids_114_0;
  reg                 ICachePlugin_logic_storage_valids_114_1;
  reg                 ICachePlugin_logic_storage_valids_115_0;
  reg                 ICachePlugin_logic_storage_valids_115_1;
  reg                 ICachePlugin_logic_storage_valids_116_0;
  reg                 ICachePlugin_logic_storage_valids_116_1;
  reg                 ICachePlugin_logic_storage_valids_117_0;
  reg                 ICachePlugin_logic_storage_valids_117_1;
  reg                 ICachePlugin_logic_storage_valids_118_0;
  reg                 ICachePlugin_logic_storage_valids_118_1;
  reg                 ICachePlugin_logic_storage_valids_119_0;
  reg                 ICachePlugin_logic_storage_valids_119_1;
  reg                 ICachePlugin_logic_storage_valids_120_0;
  reg                 ICachePlugin_logic_storage_valids_120_1;
  reg                 ICachePlugin_logic_storage_valids_121_0;
  reg                 ICachePlugin_logic_storage_valids_121_1;
  reg                 ICachePlugin_logic_storage_valids_122_0;
  reg                 ICachePlugin_logic_storage_valids_122_1;
  reg                 ICachePlugin_logic_storage_valids_123_0;
  reg                 ICachePlugin_logic_storage_valids_123_1;
  reg                 ICachePlugin_logic_storage_valids_124_0;
  reg                 ICachePlugin_logic_storage_valids_124_1;
  reg                 ICachePlugin_logic_storage_valids_125_0;
  reg                 ICachePlugin_logic_storage_valids_125_1;
  reg                 ICachePlugin_logic_storage_valids_126_0;
  reg                 ICachePlugin_logic_storage_valids_126_1;
  reg                 ICachePlugin_logic_storage_valids_127_0;
  reg                 ICachePlugin_logic_storage_valids_127_1;
  reg                 ICachePlugin_logic_tag_write_logic_fsmIsCommitting;
  reg                 ICachePlugin_logic_tag_write_logic_f2IsUpdatingLru;
  reg        [6:0]    ICachePlugin_logic_tag_write_logic_writeAddress;
  reg        [20:0]   ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag;
  reg        [20:0]   ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag;
  reg                 ICachePlugin_logic_tag_write_logic_writeData_lru;
  wire                ICachePlugin_logic_tag_write_logic_writeEnable;
  wire                ICache_F1_Access_valid;
  reg                 ICache_F2_HitCheck_valid;
  wire       [6:0]    ICachePlugin_logic_pipeline_f1_f1_index;
  wire                ICache_F1_Access_isFiring;
  wire       [20:0]   ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag;
  wire       [20:0]   ICachePlugin_logic_pipeline_f1_metaReadData_ways_1_tag;
  wire                ICachePlugin_logic_pipeline_f1_metaReadData_lru;
  wire       [42:0]   _zz_ICachePlugin_logic_pipeline_f1_metaReadData_lru;
  wire       [41:0]   _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag;
  wire       [31:0]   ICachePlugin_logic_pipeline_f1_dataReadData_0_0;
  wire       [31:0]   ICachePlugin_logic_pipeline_f1_dataReadData_0_1;
  wire       [31:0]   ICachePlugin_logic_pipeline_f1_dataReadData_0_2;
  wire       [31:0]   ICachePlugin_logic_pipeline_f1_dataReadData_0_3;
  wire       [127:0]  _zz_ICachePlugin_logic_pipeline_f1_dataReadData_0_0;
  wire       [31:0]   ICachePlugin_logic_pipeline_f1_dataReadData_1_0;
  wire       [31:0]   ICachePlugin_logic_pipeline_f1_dataReadData_1_1;
  wire       [31:0]   ICachePlugin_logic_pipeline_f1_dataReadData_1_2;
  wire       [31:0]   ICachePlugin_logic_pipeline_f1_dataReadData_1_3;
  wire       [127:0]  _zz_ICachePlugin_logic_pipeline_f1_dataReadData_1_0;
  wire                ICachePlugin_logic_pipeline_f1_writeReadHazard;
  wire       [6:0]    ICachePlugin_logic_pipeline_f2_f2_index;
  wire       [20:0]   ICachePlugin_logic_pipeline_f2_f2_tag;
  wire       [20:0]   ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_0_tag;
  wire       [20:0]   ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_1_tag;
  wire                ICachePlugin_logic_pipeline_f2_f2_metaLine_lru;
  wire                ICachePlugin_logic_pipeline_f2_hit_ways_0;
  wire                ICachePlugin_logic_pipeline_f2_hit_ways_1;
  wire                ICachePlugin_logic_pipeline_f2_isHit;
  wire       [31:0]   ICachePlugin_logic_pipeline_f2_hitWayData_0;
  wire       [31:0]   ICachePlugin_logic_pipeline_f2_hitWayData_1;
  wire       [31:0]   ICachePlugin_logic_pipeline_f2_hitWayData_2;
  wire       [31:0]   ICachePlugin_logic_pipeline_f2_hitWayData_3;
  wire                _zz_ICachePlugin_logic_pipeline_f2_hitWayIdx;
  wire       [0:0]    ICachePlugin_logic_pipeline_f2_hitWayIdx;
  wire                ICache_F2_HitCheck_isFiring;
  wire                ICachePlugin_logic_pipeline_f2_f2_can_update_lru;
  reg        [31:0]   ICachePlugin_logic_refill_refillCmdReg_address;
  reg        [7:0]    ICachePlugin_logic_refill_refillCmdReg_transactionId;
  reg        [0:0]    ICachePlugin_logic_refill_victimWayReg;
  reg        [31:0]   ICachePlugin_logic_refill_lineBuffer_0;
  reg        [31:0]   ICachePlugin_logic_refill_lineBuffer_1;
  reg        [31:0]   ICachePlugin_logic_refill_lineBuffer_2;
  reg        [31:0]   ICachePlugin_logic_refill_lineBuffer_3;
  reg                 ICachePlugin_logic_refill_refillCounter_willIncrement;
  reg                 ICachePlugin_logic_refill_refillCounter_willClear;
  reg        [1:0]    ICachePlugin_logic_refill_refillCounter_valueNext;
  reg        [1:0]    ICachePlugin_logic_refill_refillCounter_value;
  wire                ICachePlugin_logic_refill_refillCounter_willOverflowIfInc;
  wire                ICachePlugin_logic_refill_refillCounter_willOverflow;
  reg        [20:0]   ICachePlugin_logic_refill_latchedMetaOnMiss_ways_0_tag;
  reg        [20:0]   ICachePlugin_logic_refill_latchedMetaOnMiss_ways_1_tag;
  reg                 ICachePlugin_logic_refill_latchedMetaOnMiss_lru;
  wire                ICachePlugin_logic_refill_fsm_wantExit;
  reg                 ICachePlugin_logic_refill_fsm_wantStart;
  wire                ICachePlugin_logic_refill_fsm_wantKill;
  reg        [4:0]    ICachePlugin_logic_refill_fsm_stateReg;
  reg        [4:0]    ICachePlugin_logic_refill_fsm_stateNext;
  wire                when_ICachePlugin_l212;
  wire                ICachePlugin_axiMaster_ar_fire;
  wire                ICachePlugin_axiMaster_r_fire;
  wire       [3:0]    _zz_78;
  wire       [6:0]    _zz_ICachePlugin_logic_tag_write_logic_writeAddress;
  wire                when_ICachePlugin_l260;
  wire                when_ICachePlugin_l260_1;
  reg        [20:0]   _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag;
  reg        [20:0]   _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag;
  wire       [1:0]    _zz_79;
  wire       [20:0]   _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag_1;
  wire       [127:0]  _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire                _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire                _zz_152;
  wire                _zz_153;
  wire                _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire                _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire                _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire                _zz_170;
  wire                _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire                _zz_174;
  wire                _zz_175;
  wire                _zz_176;
  wire                _zz_177;
  wire                _zz_178;
  wire                _zz_179;
  wire                _zz_180;
  wire                _zz_181;
  wire                _zz_182;
  wire                _zz_183;
  wire                _zz_184;
  wire                _zz_185;
  wire                _zz_186;
  wire                _zz_187;
  wire                _zz_188;
  wire                _zz_189;
  wire                _zz_190;
  wire                _zz_191;
  wire                _zz_192;
  wire                _zz_193;
  wire                _zz_194;
  wire                _zz_195;
  wire                _zz_196;
  wire                _zz_197;
  wire                _zz_198;
  wire                _zz_199;
  wire                _zz_200;
  wire                _zz_201;
  wire                _zz_202;
  wire                _zz_203;
  wire                _zz_204;
  wire                _zz_205;
  wire                _zz_206;
  wire                _zz_207;
  wire                _zz_208;
  wire       [1:0]    _zz_209;
  wire                ICachePlugin_logic_refill_fsm_onExit_BOOT;
  wire                ICachePlugin_logic_refill_fsm_onExit_IDLE;
  wire                ICachePlugin_logic_refill_fsm_onExit_SEND_REQ;
  wire                ICachePlugin_logic_refill_fsm_onExit_RECEIVE_DATA;
  wire                ICachePlugin_logic_refill_fsm_onExit_COMMIT;
  wire                ICachePlugin_logic_refill_fsm_onEntry_BOOT;
  wire                ICachePlugin_logic_refill_fsm_onEntry_IDLE;
  wire                ICachePlugin_logic_refill_fsm_onEntry_SEND_REQ;
  wire                ICachePlugin_logic_refill_fsm_onEntry_RECEIVE_DATA;
  wire                ICachePlugin_logic_refill_fsm_onEntry_COMMIT;
  reg        [2:0]    ICachePlugin_logic_management_sim_fsmStateId;
  wire                when_ICachePlugin_l299;
  wire                when_ICachePlugin_l300;
  wire                when_ICachePlugin_l301;
  wire                when_ICachePlugin_l302;
  wire                BpuPipelinePlugin_logic_s1_read_valid;
  reg                 BpuPipelinePlugin_logic_s2_predict_valid;
  wire                BpuPipelinePlugin_logic_s1_read_isFiring;
  wire       [9:0]    _zz_210;
  wire       [7:0]    _zz_211;
  wire       [9:0]    _zz_BpuPipelinePlugin_logic_phtReadData_s1;
  wire       [1:0]    BpuPipelinePlugin_logic_phtReadData_s1;
  wire       [7:0]    _zz_BpuPipelinePlugin_logic_btbReadData_s1_valid;
  wire                BpuPipelinePlugin_logic_btbReadData_s1_valid;
  wire       [21:0]   BpuPipelinePlugin_logic_btbReadData_s1_tag;
  wire       [31:0]   BpuPipelinePlugin_logic_btbReadData_s1_target;
  wire       [54:0]   _zz_BpuPipelinePlugin_logic_btbReadData_s1_valid_1;
  wire                BpuPipelinePlugin_logic_phtPrediction;
  wire                BpuPipelinePlugin_logic_btbHit;
  wire                BpuPipelinePlugin_logic_s2_predict_isFiring;
  wire                _zz_214;
  wire                BpuPipelinePlugin_logic_u1_read_valid;
  reg                 BpuPipelinePlugin_logic_u2_write_valid;
  wire                BpuPipelinePlugin_logic_u1_read_isFiring;
  wire       [9:0]    _zz_BpuPipelinePlugin_logic_oldPhtState_u1;
  wire       [1:0]    BpuPipelinePlugin_logic_oldPhtState_u1;
  reg        [1:0]    BpuPipelinePlugin_logic_newPhtState;
  wire                BpuPipelinePlugin_logic_u2_write_isFiring;
  reg        [31:0]   BpuPipelinePlugin_queryPortIn_payload_pc_regNext;
  reg        [2:0]    BpuPipelinePlugin_queryPortIn_payload_transactionId_regNext;
  wire                uartAxi_aw_valid;
  wire                uartAxi_aw_ready;
  wire       [31:0]   uartAxi_aw_payload_addr;
  wire       [6:0]    uartAxi_aw_payload_id;
  wire       [7:0]    uartAxi_aw_payload_len;
  wire       [2:0]    uartAxi_aw_payload_size;
  wire       [1:0]    uartAxi_aw_payload_burst;
  wire                uartAxi_w_valid;
  wire                uartAxi_w_ready;
  wire       [31:0]   uartAxi_w_payload_data;
  wire       [3:0]    uartAxi_w_payload_strb;
  wire                uartAxi_w_payload_last;
  wire                uartAxi_b_valid;
  wire                uartAxi_b_ready;
  wire       [6:0]    uartAxi_b_payload_id;
  wire       [1:0]    uartAxi_b_payload_resp;
  wire                uartAxi_ar_valid;
  wire                uartAxi_ar_ready;
  wire       [31:0]   uartAxi_ar_payload_addr;
  wire       [6:0]    uartAxi_ar_payload_id;
  wire       [7:0]    uartAxi_ar_payload_len;
  wire       [2:0]    uartAxi_ar_payload_size;
  wire       [1:0]    uartAxi_ar_payload_burst;
  wire                uartAxi_r_valid;
  wire                uartAxi_r_ready;
  wire       [31:0]   uartAxi_r_payload_data;
  wire       [6:0]    uartAxi_r_payload_id;
  wire       [1:0]    uartAxi_r_payload_resp;
  wire                uartAxi_r_payload_last;
  wire                io_axiOut_readOnly_ar_valid;
  wire                io_axiOut_readOnly_ar_ready;
  wire       [31:0]   io_axiOut_readOnly_ar_payload_addr;
  wire       [3:0]    io_axiOut_readOnly_ar_payload_id;
  wire       [7:0]    io_axiOut_readOnly_ar_payload_len;
  wire       [2:0]    io_axiOut_readOnly_ar_payload_size;
  wire       [1:0]    io_axiOut_readOnly_ar_payload_burst;
  wire                io_axiOut_readOnly_r_valid;
  wire                io_axiOut_readOnly_r_ready;
  wire       [31:0]   io_axiOut_readOnly_r_payload_data;
  wire       [3:0]    io_axiOut_readOnly_r_payload_id;
  wire       [1:0]    io_axiOut_readOnly_r_payload_resp;
  wire                io_axiOut_readOnly_r_payload_last;
  wire                io_axiOut_writeOnly_aw_valid;
  wire                io_axiOut_writeOnly_aw_ready;
  wire       [31:0]   io_axiOut_writeOnly_aw_payload_addr;
  wire       [3:0]    io_axiOut_writeOnly_aw_payload_id;
  wire       [7:0]    io_axiOut_writeOnly_aw_payload_len;
  wire       [2:0]    io_axiOut_writeOnly_aw_payload_size;
  wire       [1:0]    io_axiOut_writeOnly_aw_payload_burst;
  wire                io_axiOut_writeOnly_w_valid;
  wire                io_axiOut_writeOnly_w_ready;
  wire       [31:0]   io_axiOut_writeOnly_w_payload_data;
  wire       [3:0]    io_axiOut_writeOnly_w_payload_strb;
  wire                io_axiOut_writeOnly_w_payload_last;
  wire                io_axiOut_writeOnly_b_valid;
  wire                io_axiOut_writeOnly_b_ready;
  wire       [3:0]    io_axiOut_writeOnly_b_payload_id;
  wire       [1:0]    io_axiOut_writeOnly_b_payload_resp;
  wire                io_axiOut_readOnly_ar_valid_1;
  wire                io_axiOut_readOnly_ar_ready_1;
  wire       [31:0]   io_axiOut_readOnly_ar_payload_addr_1;
  wire       [3:0]    io_axiOut_readOnly_ar_payload_id_1;
  wire       [7:0]    io_axiOut_readOnly_ar_payload_len_1;
  wire       [2:0]    io_axiOut_readOnly_ar_payload_size_1;
  wire       [1:0]    io_axiOut_readOnly_ar_payload_burst_1;
  wire                io_axiOut_readOnly_r_valid_1;
  wire                io_axiOut_readOnly_r_ready_1;
  wire       [31:0]   io_axiOut_readOnly_r_payload_data_1;
  wire       [3:0]    io_axiOut_readOnly_r_payload_id_1;
  wire       [1:0]    io_axiOut_readOnly_r_payload_resp_1;
  wire                io_axiOut_readOnly_r_payload_last_1;
  wire                io_axiOut_writeOnly_aw_valid_1;
  wire                io_axiOut_writeOnly_aw_ready_1;
  wire       [31:0]   io_axiOut_writeOnly_aw_payload_addr_1;
  wire       [3:0]    io_axiOut_writeOnly_aw_payload_id_1;
  wire       [7:0]    io_axiOut_writeOnly_aw_payload_len_1;
  wire       [2:0]    io_axiOut_writeOnly_aw_payload_size_1;
  wire       [1:0]    io_axiOut_writeOnly_aw_payload_burst_1;
  wire                io_axiOut_writeOnly_w_valid_1;
  wire                io_axiOut_writeOnly_w_ready_1;
  wire       [31:0]   io_axiOut_writeOnly_w_payload_data_1;
  wire       [3:0]    io_axiOut_writeOnly_w_payload_strb_1;
  wire                io_axiOut_writeOnly_w_payload_last_1;
  wire                io_axiOut_writeOnly_b_valid_1;
  wire                io_axiOut_writeOnly_b_ready_1;
  wire       [3:0]    io_axiOut_writeOnly_b_payload_id_1;
  wire       [1:0]    io_axiOut_writeOnly_b_payload_resp_1;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_ar_valid;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_ar_ready;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_r_valid;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_r_ready;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_data;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_id;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_resp;
  wire                DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_last;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_aw_valid;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_aw_ready;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_addr;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_id;
  wire       [7:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_len;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_size;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_burst;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_prot;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_w_valid;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_w_ready;
  wire       [31:0]   DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_data;
  wire       [3:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_strb;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_last;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_b_valid;
  wire                DataCachePlugin_setup_dcacheMaster_writeOnly_b_ready;
  wire       [2:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_b_payload_id;
  wire       [1:0]    DataCachePlugin_setup_dcacheMaster_writeOnly_b_payload_resp;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_ready;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_r_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_r_ready;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_id;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_resp;
  wire                CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_last;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_ready;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_addr;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_id;
  wire       [7:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_len;
  wire       [2:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_size;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_burst;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_ready;
  wire       [31:0]   CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_data;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_strb;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_last;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_valid;
  wire                CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_ready;
  wire       [3:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_payload_id;
  wire       [1:0]    CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_payload_resp;
  wire                io_outputs_0_ar_validPipe_valid;
  wire                io_outputs_0_ar_validPipe_ready;
  wire       [31:0]   io_outputs_0_ar_validPipe_payload_addr;
  wire       [3:0]    io_outputs_0_ar_validPipe_payload_id;
  wire       [7:0]    io_outputs_0_ar_validPipe_payload_len;
  wire       [2:0]    io_outputs_0_ar_validPipe_payload_size;
  wire       [1:0]    io_outputs_0_ar_validPipe_payload_burst;
  reg                 io_outputs_0_ar_rValid;
  wire                io_outputs_0_ar_validPipe_fire;
  wire                io_outputs_1_ar_validPipe_valid;
  wire                io_outputs_1_ar_validPipe_ready;
  wire       [31:0]   io_outputs_1_ar_validPipe_payload_addr;
  wire       [3:0]    io_outputs_1_ar_validPipe_payload_id;
  wire       [7:0]    io_outputs_1_ar_validPipe_payload_len;
  wire       [2:0]    io_outputs_1_ar_validPipe_payload_size;
  wire       [1:0]    io_outputs_1_ar_validPipe_payload_burst;
  reg                 io_outputs_1_ar_rValid;
  wire                io_outputs_1_ar_validPipe_fire;
  wire                io_outputs_2_ar_validPipe_valid;
  wire                io_outputs_2_ar_validPipe_ready;
  wire       [31:0]   io_outputs_2_ar_validPipe_payload_addr;
  wire       [3:0]    io_outputs_2_ar_validPipe_payload_id;
  wire       [7:0]    io_outputs_2_ar_validPipe_payload_len;
  wire       [2:0]    io_outputs_2_ar_validPipe_payload_size;
  wire       [1:0]    io_outputs_2_ar_validPipe_payload_burst;
  reg                 io_outputs_2_ar_rValid;
  wire                io_outputs_2_ar_validPipe_fire;
  wire                io_outputs_0_aw_validPipe_valid;
  wire                io_outputs_0_aw_validPipe_ready;
  wire       [31:0]   io_outputs_0_aw_validPipe_payload_addr;
  wire       [3:0]    io_outputs_0_aw_validPipe_payload_id;
  wire       [7:0]    io_outputs_0_aw_validPipe_payload_len;
  wire       [2:0]    io_outputs_0_aw_validPipe_payload_size;
  wire       [1:0]    io_outputs_0_aw_validPipe_payload_burst;
  reg                 io_outputs_0_aw_rValid;
  wire                io_outputs_0_aw_validPipe_fire;
  wire                io_outputs_1_aw_validPipe_valid;
  wire                io_outputs_1_aw_validPipe_ready;
  wire       [31:0]   io_outputs_1_aw_validPipe_payload_addr;
  wire       [3:0]    io_outputs_1_aw_validPipe_payload_id;
  wire       [7:0]    io_outputs_1_aw_validPipe_payload_len;
  wire       [2:0]    io_outputs_1_aw_validPipe_payload_size;
  wire       [1:0]    io_outputs_1_aw_validPipe_payload_burst;
  reg                 io_outputs_1_aw_rValid;
  wire                io_outputs_1_aw_validPipe_fire;
  wire                io_outputs_2_aw_validPipe_valid;
  wire                io_outputs_2_aw_validPipe_ready;
  wire       [31:0]   io_outputs_2_aw_validPipe_payload_addr;
  wire       [3:0]    io_outputs_2_aw_validPipe_payload_id;
  wire       [7:0]    io_outputs_2_aw_validPipe_payload_len;
  wire       [2:0]    io_outputs_2_aw_validPipe_payload_size;
  wire       [1:0]    io_outputs_2_aw_validPipe_payload_burst;
  reg                 io_outputs_2_aw_rValid;
  wire                io_outputs_2_aw_validPipe_fire;
  wire                io_outputs_0_ar_validPipe_valid_1;
  wire                io_outputs_0_ar_validPipe_ready_1;
  wire       [31:0]   io_outputs_0_ar_validPipe_payload_addr_1;
  wire       [3:0]    io_outputs_0_ar_validPipe_payload_id_1;
  wire       [7:0]    io_outputs_0_ar_validPipe_payload_len_1;
  wire       [2:0]    io_outputs_0_ar_validPipe_payload_size_1;
  wire       [1:0]    io_outputs_0_ar_validPipe_payload_burst_1;
  reg                 io_outputs_0_ar_rValid_1;
  wire                io_outputs_0_ar_validPipe_fire_1;
  wire                io_outputs_1_ar_validPipe_valid_1;
  wire                io_outputs_1_ar_validPipe_ready_1;
  wire       [31:0]   io_outputs_1_ar_validPipe_payload_addr_1;
  wire       [3:0]    io_outputs_1_ar_validPipe_payload_id_1;
  wire       [7:0]    io_outputs_1_ar_validPipe_payload_len_1;
  wire       [2:0]    io_outputs_1_ar_validPipe_payload_size_1;
  wire       [1:0]    io_outputs_1_ar_validPipe_payload_burst_1;
  reg                 io_outputs_1_ar_rValid_1;
  wire                io_outputs_1_ar_validPipe_fire_1;
  wire                io_outputs_2_ar_validPipe_valid_1;
  wire                io_outputs_2_ar_validPipe_ready_1;
  wire       [31:0]   io_outputs_2_ar_validPipe_payload_addr_1;
  wire       [3:0]    io_outputs_2_ar_validPipe_payload_id_1;
  wire       [7:0]    io_outputs_2_ar_validPipe_payload_len_1;
  wire       [2:0]    io_outputs_2_ar_validPipe_payload_size_1;
  wire       [1:0]    io_outputs_2_ar_validPipe_payload_burst_1;
  reg                 io_outputs_2_ar_rValid_1;
  wire                io_outputs_2_ar_validPipe_fire_1;
  wire                io_outputs_0_aw_validPipe_valid_1;
  wire                io_outputs_0_aw_validPipe_ready_1;
  wire       [31:0]   io_outputs_0_aw_validPipe_payload_addr_1;
  wire       [3:0]    io_outputs_0_aw_validPipe_payload_id_1;
  wire       [7:0]    io_outputs_0_aw_validPipe_payload_len_1;
  wire       [2:0]    io_outputs_0_aw_validPipe_payload_size_1;
  wire       [1:0]    io_outputs_0_aw_validPipe_payload_burst_1;
  reg                 io_outputs_0_aw_rValid_1;
  wire                io_outputs_0_aw_validPipe_fire_1;
  wire                io_outputs_1_aw_validPipe_valid_1;
  wire                io_outputs_1_aw_validPipe_ready_1;
  wire       [31:0]   io_outputs_1_aw_validPipe_payload_addr_1;
  wire       [3:0]    io_outputs_1_aw_validPipe_payload_id_1;
  wire       [7:0]    io_outputs_1_aw_validPipe_payload_len_1;
  wire       [2:0]    io_outputs_1_aw_validPipe_payload_size_1;
  wire       [1:0]    io_outputs_1_aw_validPipe_payload_burst_1;
  reg                 io_outputs_1_aw_rValid_1;
  wire                io_outputs_1_aw_validPipe_fire_1;
  wire                io_outputs_2_aw_validPipe_valid_1;
  wire                io_outputs_2_aw_validPipe_ready_1;
  wire       [31:0]   io_outputs_2_aw_validPipe_payload_addr_1;
  wire       [3:0]    io_outputs_2_aw_validPipe_payload_id_1;
  wire       [7:0]    io_outputs_2_aw_validPipe_payload_len_1;
  wire       [2:0]    io_outputs_2_aw_validPipe_payload_size_1;
  wire       [1:0]    io_outputs_2_aw_validPipe_payload_burst_1;
  reg                 io_outputs_2_aw_rValid_1;
  wire                io_outputs_2_aw_validPipe_fire_1;
  wire                io_outputs_0_ar_validPipe_valid_2;
  wire                io_outputs_0_ar_validPipe_ready_2;
  wire       [31:0]   io_outputs_0_ar_validPipe_payload_addr_2;
  wire       [2:0]    io_outputs_0_ar_validPipe_payload_id_2;
  wire       [7:0]    io_outputs_0_ar_validPipe_payload_len_2;
  wire       [2:0]    io_outputs_0_ar_validPipe_payload_size_2;
  wire       [1:0]    io_outputs_0_ar_validPipe_payload_burst_2;
  wire       [2:0]    io_outputs_0_ar_validPipe_payload_prot;
  reg                 io_outputs_0_ar_rValid_2;
  wire                io_outputs_0_ar_validPipe_fire_2;
  wire                io_outputs_1_ar_validPipe_valid_2;
  wire                io_outputs_1_ar_validPipe_ready_2;
  wire       [31:0]   io_outputs_1_ar_validPipe_payload_addr_2;
  wire       [2:0]    io_outputs_1_ar_validPipe_payload_id_2;
  wire       [7:0]    io_outputs_1_ar_validPipe_payload_len_2;
  wire       [2:0]    io_outputs_1_ar_validPipe_payload_size_2;
  wire       [1:0]    io_outputs_1_ar_validPipe_payload_burst_2;
  wire       [2:0]    io_outputs_1_ar_validPipe_payload_prot;
  reg                 io_outputs_1_ar_rValid_2;
  wire                io_outputs_1_ar_validPipe_fire_2;
  wire                io_outputs_2_ar_validPipe_valid_2;
  wire                io_outputs_2_ar_validPipe_ready_2;
  wire       [31:0]   io_outputs_2_ar_validPipe_payload_addr_2;
  wire       [2:0]    io_outputs_2_ar_validPipe_payload_id_2;
  wire       [7:0]    io_outputs_2_ar_validPipe_payload_len_2;
  wire       [2:0]    io_outputs_2_ar_validPipe_payload_size_2;
  wire       [1:0]    io_outputs_2_ar_validPipe_payload_burst_2;
  wire       [2:0]    io_outputs_2_ar_validPipe_payload_prot;
  reg                 io_outputs_2_ar_rValid_2;
  wire                io_outputs_2_ar_validPipe_fire_2;
  wire                io_outputs_0_aw_validPipe_valid_2;
  wire                io_outputs_0_aw_validPipe_ready_2;
  wire       [31:0]   io_outputs_0_aw_validPipe_payload_addr_2;
  wire       [2:0]    io_outputs_0_aw_validPipe_payload_id_2;
  wire       [7:0]    io_outputs_0_aw_validPipe_payload_len_2;
  wire       [2:0]    io_outputs_0_aw_validPipe_payload_size_2;
  wire       [1:0]    io_outputs_0_aw_validPipe_payload_burst_2;
  wire       [2:0]    io_outputs_0_aw_validPipe_payload_prot;
  reg                 io_outputs_0_aw_rValid_2;
  wire                io_outputs_0_aw_validPipe_fire_2;
  wire                io_outputs_1_aw_validPipe_valid_2;
  wire                io_outputs_1_aw_validPipe_ready_2;
  wire       [31:0]   io_outputs_1_aw_validPipe_payload_addr_2;
  wire       [2:0]    io_outputs_1_aw_validPipe_payload_id_2;
  wire       [7:0]    io_outputs_1_aw_validPipe_payload_len_2;
  wire       [2:0]    io_outputs_1_aw_validPipe_payload_size_2;
  wire       [1:0]    io_outputs_1_aw_validPipe_payload_burst_2;
  wire       [2:0]    io_outputs_1_aw_validPipe_payload_prot;
  reg                 io_outputs_1_aw_rValid_2;
  wire                io_outputs_1_aw_validPipe_fire_2;
  wire                io_outputs_2_aw_validPipe_valid_2;
  wire                io_outputs_2_aw_validPipe_ready_2;
  wire       [31:0]   io_outputs_2_aw_validPipe_payload_addr_2;
  wire       [2:0]    io_outputs_2_aw_validPipe_payload_id_2;
  wire       [7:0]    io_outputs_2_aw_validPipe_payload_len_2;
  wire       [2:0]    io_outputs_2_aw_validPipe_payload_size_2;
  wire       [1:0]    io_outputs_2_aw_validPipe_payload_burst_2;
  wire       [2:0]    io_outputs_2_aw_validPipe_payload_prot;
  reg                 io_outputs_2_aw_rValid_2;
  wire                io_outputs_2_aw_validPipe_fire_2;
  wire                io_outputs_0_ar_validPipe_valid_3;
  wire                io_outputs_0_ar_validPipe_ready_3;
  wire       [31:0]   io_outputs_0_ar_validPipe_payload_addr_3;
  wire       [3:0]    io_outputs_0_ar_validPipe_payload_id_3;
  wire       [7:0]    io_outputs_0_ar_validPipe_payload_len_3;
  wire       [2:0]    io_outputs_0_ar_validPipe_payload_size_3;
  wire       [1:0]    io_outputs_0_ar_validPipe_payload_burst_3;
  reg                 io_outputs_0_ar_rValid_3;
  wire                io_outputs_0_ar_validPipe_fire_3;
  wire                io_outputs_1_ar_validPipe_valid_3;
  wire                io_outputs_1_ar_validPipe_ready_3;
  wire       [31:0]   io_outputs_1_ar_validPipe_payload_addr_3;
  wire       [3:0]    io_outputs_1_ar_validPipe_payload_id_3;
  wire       [7:0]    io_outputs_1_ar_validPipe_payload_len_3;
  wire       [2:0]    io_outputs_1_ar_validPipe_payload_size_3;
  wire       [1:0]    io_outputs_1_ar_validPipe_payload_burst_3;
  reg                 io_outputs_1_ar_rValid_3;
  wire                io_outputs_1_ar_validPipe_fire_3;
  wire                io_outputs_2_ar_validPipe_valid_3;
  wire                io_outputs_2_ar_validPipe_ready_3;
  wire       [31:0]   io_outputs_2_ar_validPipe_payload_addr_3;
  wire       [3:0]    io_outputs_2_ar_validPipe_payload_id_3;
  wire       [7:0]    io_outputs_2_ar_validPipe_payload_len_3;
  wire       [2:0]    io_outputs_2_ar_validPipe_payload_size_3;
  wire       [1:0]    io_outputs_2_ar_validPipe_payload_burst_3;
  reg                 io_outputs_2_ar_rValid_3;
  wire                io_outputs_2_ar_validPipe_fire_3;
  wire                io_outputs_0_aw_validPipe_valid_3;
  wire                io_outputs_0_aw_validPipe_ready_3;
  wire       [31:0]   io_outputs_0_aw_validPipe_payload_addr_3;
  wire       [3:0]    io_outputs_0_aw_validPipe_payload_id_3;
  wire       [7:0]    io_outputs_0_aw_validPipe_payload_len_3;
  wire       [2:0]    io_outputs_0_aw_validPipe_payload_size_3;
  wire       [1:0]    io_outputs_0_aw_validPipe_payload_burst_3;
  reg                 io_outputs_0_aw_rValid_3;
  wire                io_outputs_0_aw_validPipe_fire_3;
  wire                io_outputs_1_aw_validPipe_valid_3;
  wire                io_outputs_1_aw_validPipe_ready_3;
  wire       [31:0]   io_outputs_1_aw_validPipe_payload_addr_3;
  wire       [3:0]    io_outputs_1_aw_validPipe_payload_id_3;
  wire       [7:0]    io_outputs_1_aw_validPipe_payload_len_3;
  wire       [2:0]    io_outputs_1_aw_validPipe_payload_size_3;
  wire       [1:0]    io_outputs_1_aw_validPipe_payload_burst_3;
  reg                 io_outputs_1_aw_rValid_3;
  wire                io_outputs_1_aw_validPipe_fire_3;
  wire                io_outputs_2_aw_validPipe_valid_3;
  wire                io_outputs_2_aw_validPipe_ready_3;
  wire       [31:0]   io_outputs_2_aw_validPipe_payload_addr_3;
  wire       [3:0]    io_outputs_2_aw_validPipe_payload_id_3;
  wire       [7:0]    io_outputs_2_aw_validPipe_payload_len_3;
  wire       [2:0]    io_outputs_2_aw_validPipe_payload_size_3;
  wire       [1:0]    io_outputs_2_aw_validPipe_payload_burst_3;
  reg                 io_outputs_2_aw_rValid_3;
  wire                io_outputs_2_aw_validPipe_fire_3;
  reg                 _zz_io_leds;
  wire                _zz_when_CoreNSCSCC_l598;
  reg                 _zz_when_CoreNSCSCC_l598_1;
  wire                when_CoreNSCSCC_l598;
  `ifndef SYNTHESIS
  reg [87:0] _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string;
  reg [39:0] _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string;
  reg [87:0] _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string;
  reg [39:0] _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1_string;
  reg [87:0] _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string;
  reg [39:0] _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2_string;
  reg [87:0] _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string;
  reg [39:0] _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3_string;
  reg [127:0] _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_string;
  reg [39:0] _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string;
  reg [103:0] _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string;
  reg [127:0] _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_1_string;
  reg [39:0] _zz_io_iqEntryIn_payload_aluCtrl_logicOp_string;
  reg [103:0] _zz_io_iqEntryIn_payload_immUsage_string;
  reg [39:0] _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1_string;
  reg [103:0] _zz_io_iqEntryIn_payload_immUsage_1_string;
  reg [39:0] _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2_string;
  reg [103:0] _zz_io_iqEntryIn_payload_immUsage_2_string;
  reg [87:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string;
  reg [151:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string;
  reg [71:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string;
  reg [103:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string;
  reg [87:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string;
  reg [87:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string;
  reg [151:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string;
  reg [71:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype_string;
  reg [103:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size_string;
  reg [87:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode_string;
  reg [87:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string;
  reg [151:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string;
  reg [71:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string;
  reg [103:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string;
  reg [87:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string;
  reg [39:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string;
  reg [95:0] s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string;
  reg [87:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string;
  reg [151:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string;
  reg [71:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa_string;
  reg [39:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string;
  reg [39:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string;
  reg [39:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string;
  reg [103:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string;
  reg [39:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string;
  reg [7:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string;
  reg [87:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string;
  reg [39:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string;
  reg [7:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string;
  reg [95:0] s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string;
  reg [87:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string;
  reg [151:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string;
  reg [71:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string;
  reg [39:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string;
  reg [39:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string;
  reg [39:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string;
  reg [103:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string;
  reg [39:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string;
  reg [7:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string;
  reg [87:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string;
  reg [39:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string;
  reg [87:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string;
  reg [151:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string;
  reg [71:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa_string;
  reg [39:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string;
  reg [39:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string;
  reg [39:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string;
  reg [103:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string;
  reg [39:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string;
  reg [7:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string;
  reg [87:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string;
  reg [39:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string;
  reg [7:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string;
  reg [95:0] s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string;
  reg [151:0] ROBPlugin_aggregatedFlushSignal_payload_reason_string;
  reg [39:0] AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string;
  reg [103:0] AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_0_0_0_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_0_0_1_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_0_0_2_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_0_0_3_string;
  reg [87:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string;
  reg [151:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string;
  reg [71:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa_string;
  reg [39:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype_string;
  reg [39:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype_string;
  reg [39:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype_string;
  reg [103:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string;
  reg [39:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size_string;
  reg [87:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string;
  reg [39:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_1_0_0_string;
  reg [87:0] BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string;
  reg [39:0] BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_2_0_0_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_2_0_1_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_2_0_2_string;
  reg [7:0] LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_3_0_0_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_3_0_1_string;
  reg [151:0] CommitPlugin_hw_robFlushPort_payload_reason_string;
  reg [7:0] LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize_string;
  reg [7:0] LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string;
  reg [7:0] StoreBufferPlugin_hw_pushPortInst_payload_accessSize_string;
  reg [7:0] StoreBufferPlugin_hw_bypassQuerySizeIn_string;
  reg [7:0] StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size_string;
  reg [7:0] LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size_string;
  reg [87:0] DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string;
  reg [151:0] DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string;
  reg [71:0] DecodePlugin_logic_decodedUopsOutputVec_0_isa_string;
  reg [39:0] DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string;
  reg [39:0] DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string;
  reg [39:0] DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string;
  reg [103:0] DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string;
  reg [39:0] DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string;
  reg [7:0] DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string;
  reg [87:0] DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string;
  reg [39:0] DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string;
  reg [7:0] DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string;
  reg [95:0] DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string;
  reg [87:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string;
  reg [151:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string;
  reg [71:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa_string;
  reg [39:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string;
  reg [39:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string;
  reg [39:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string;
  reg [103:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string;
  reg [39:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string;
  reg [7:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string;
  reg [87:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string;
  reg [39:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string;
  reg [7:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string;
  reg [95:0] _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string;
  reg [39:0] DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype_string;
  reg [87:0] RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string;
  reg [151:0] RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string;
  reg [71:0] RobAllocPlugin_logic_allocatedUops_0_decoded_isa_string;
  reg [39:0] RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype_string;
  reg [39:0] RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype_string;
  reg [39:0] RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype_string;
  reg [103:0] RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string;
  reg [39:0] RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp_string;
  reg [7:0] RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size_string;
  reg [87:0] RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string;
  reg [39:0] RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string;
  reg [151:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string;
  reg [71:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string;
  reg [151:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string;
  reg [71:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string;
  reg [151:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string;
  reg [71:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string;
  reg [151:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string;
  reg [71:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode_string;
  reg [39:0] AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp_string;
  reg [103:0] AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string;
  reg [87:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string;
  reg [151:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string;
  reg [71:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa_string;
  reg [39:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string;
  reg [39:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string;
  reg [39:0] BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype_string;
  reg [7:0] LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size_string;
  reg [7:0] _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string;
  reg [7:0] LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string;
  reg [7:0] io_outputs_0_combStage_payload_accessSize_string;
  reg [7:0] io_outputs_1_combStage_payload_accessSize_string;
  reg [7:0] _zz_io_outputs_0_combStage_translated_payload_size_string;
  reg [7:0] io_outputs_0_combStage_translated_payload_size_string;
  reg [7:0] _zz_io_outputs_1_combStage_translated_payload_accessSize_string;
  reg [7:0] io_outputs_1_combStage_translated_payload_accessSize_string;
  reg [7:0] _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_string;
  reg [7:0] _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string;
  reg [7:0] _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1_string;
  reg [7:0] _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2_string;
  reg [7:0] LoadQueuePlugin_logic_pushCmd_payload_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slots_0_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slots_1_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slots_2_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slots_3_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slotsNext_0_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slotsNext_1_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slotsNext_2_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_slotsNext_3_size_string;
  reg [7:0] LoadQueuePlugin_logic_loadQueue_completingHead_size_string;
  reg [7:0] StoreBufferPlugin_logic_slots_0_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slots_1_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slots_2_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slots_3_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slotsNext_0_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slotsNext_1_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slotsNext_2_accessSize_string;
  reg [7:0] StoreBufferPlugin_logic_slotsNext_3_accessSize_string;
  reg [7:0] _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string;
  reg [151:0] _zz_ROBPlugin_aggregatedFlushSignal_payload_reason_string;
  reg [95:0] ICachePlugin_logic_refill_fsm_stateReg_string;
  reg [95:0] ICachePlugin_logic_refill_fsm_stateNext_string;
  `endif

  (* ram_style = "block" *) reg [42:0] ICachePlugin_logic_storage_tagLruRam [0:127];
  (* ram_style = "block" *) reg [127:0] ICachePlugin_logic_storage_dataRams_0 [0:127];
  (* ram_style = "block" *) reg [127:0] ICachePlugin_logic_storage_dataRams_1 [0:127];
  (* ram_style = "block" *) reg [1:0] BpuPipelinePlugin_logic_pht [0:1023];
  (* ram_style = "block" *) reg [54:0] BpuPipelinePlugin_logic_btb [0:255];
  function [63:0] zz_CheckpointManagerPlugin_logic_initialFreeMask(input dummy);
    begin
      zz_CheckpointManagerPlugin_logic_initialFreeMask = 64'h0;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[32] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[33] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[34] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[35] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[36] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[37] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[38] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[39] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[40] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[41] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[42] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[43] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[44] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[45] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[46] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[47] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[48] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[49] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[50] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[51] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[52] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[53] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[54] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[55] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[56] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[57] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[58] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[59] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[60] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[61] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[62] = 1'b1;
      zz_CheckpointManagerPlugin_logic_initialFreeMask[63] = 1'b1;
    end
  endfunction
  wire [63:0] _zz_220;

  assign _zz_io_triggerIn_1 = 1'b1;
  assign _zz_io_triggerIn = {7'd0, _zz_io_triggerIn_1};
  assign _zz_when_Debug_l71_13 = {7'd0, _zz_when_Debug_l71_1};
  assign _zz_io_triggerIn_3 = 5'h13;
  assign _zz_io_triggerIn_2 = {3'd0, _zz_io_triggerIn_3};
  assign _zz_when_Debug_l71_1_1 = {3'd0, _zz_when_Debug_l71_2};
  assign _zz_io_triggerIn_5 = 5'h15;
  assign _zz_io_triggerIn_4 = {3'd0, _zz_io_triggerIn_5};
  assign _zz_when_Debug_l71_2_1 = {3'd0, _zz_when_Debug_l71_3};
  assign _zz_io_triggerIn_7 = 5'h14;
  assign _zz_io_triggerIn_6 = {3'd0, _zz_io_triggerIn_7};
  assign _zz_when_Debug_l71_3_1 = {3'd0, _zz_when_Debug_l71_4};
  assign _zz_io_triggerIn_9 = 5'h16;
  assign _zz_io_triggerIn_8 = {3'd0, _zz_io_triggerIn_9};
  assign _zz_when_Debug_l71_4_1 = {3'd0, _zz_when_Debug_l71_5};
  assign _zz_CommitPlugin_commitStatsReg_totalCommitted = {31'd0, CommitPlugin_logic_s1_s1_committedThisCycle};
  assign _zz_CommitPlugin_commitStatsReg_physRegRecycled = {31'd0, CommitPlugin_logic_s1_s1_recycledThisCycle};
  assign _zz_CommitPlugin_commitStatsReg_robFlushCount = {31'd0, CommitPlugin_logic_s1_s1_flushedThisCycle};
  assign _zz_io_triggerIn_11 = 5'h19;
  assign _zz_io_triggerIn_10 = {3'd0, _zz_io_triggerIn_11};
  assign _zz_when_Debug_l71_5_1 = {3'd0, _zz_when_Debug_l71_6};
  assign _zz_io_triggerIn_13 = 5'h17;
  assign _zz_io_triggerIn_12 = {3'd0, _zz_io_triggerIn_13};
  assign _zz_when_Debug_l71_6_1 = {3'd0, _zz_when_Debug_l71_7};
  assign _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_2 = _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode;
  assign _zz_io_triggerIn_15 = 5'h18;
  assign _zz_io_triggerIn_14 = {3'd0, _zz_io_triggerIn_15};
  assign _zz_when_Debug_l71_7_1 = {3'd0, _zz_when_Debug_l71_8};
  assign _zz_MulEU_MulEuPlugin_euResult_data_1 = _zz_MulEU_MulEuPlugin_euResult_data;
  assign _zz_io_triggerIn_17 = 5'h18;
  assign _zz_io_triggerIn_16 = {3'd0, _zz_io_triggerIn_17};
  assign _zz_when_Debug_l71_8_1 = {3'd0, _zz_when_Debug_l71_9};
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3 = BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_1 = BranchEU_BranchEuPlugin_gprReadPorts_1_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_2 = BranchEU_BranchEuPlugin_gprReadPorts_1_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_3 = BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_4 = BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_5 = BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_6 = BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_7 = BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4 = _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_2;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_1 = ($signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_2) + $signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_3));
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_2 = BranchEU_BranchEuPlugin_gprReadPorts_0_rsp;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_3 = _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_2;
  assign _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_4 = _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_2;
  assign _zz_io_triggerIn_19 = 5'h18;
  assign _zz_io_triggerIn_18 = {3'd0, _zz_io_triggerIn_19};
  assign _zz_when_Debug_l71_9_1 = {3'd0, _zz_when_Debug_l71_10};
  assign _zz_io_triggerIn_21 = 5'h18;
  assign _zz_io_triggerIn_20 = {3'd0, _zz_io_triggerIn_21};
  assign _zz_when_Debug_l71_10_1 = {3'd0, _zz_when_Debug_l71_11};
  assign _zz__zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_2 = {29'd0, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_1};
  assign _zz_LoadQueuePlugin_logic_loadQueue_pushOh = ((~ LoadQueuePlugin_logic_loadQueue_availableSlotsMask) + 4'b0001);
  assign _zz_StoreBufferPlugin_logic_dcacheResponseForHead = StoreBufferPlugin_logic_slots_0_robPtr[2:0];
  assign _zz_io_triggerIn_23 = 6'h20;
  assign _zz_io_triggerIn_22 = {2'd0, _zz_io_triggerIn_23};
  assign _zz_when_Debug_l71_11_1 = {2'd0, _zz_when_Debug_l71_12};
  assign _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_1 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[1 : 0];
  assign _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask = ({3'd0,1'b1} <<< _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_1);
  assign _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_2 = _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_3;
  assign _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_3 = ({3'd0,2'b11} <<< _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_4);
  assign _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_4 = ({1'd0,_zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_1[1 : 1]} <<< 1'd1);
  assign _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_5 = _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_6;
  assign _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_6 = ({3'd0,4'b1111} <<< 2'b00);
  assign _zz__zz_StoreBufferPlugin_logic_loadQueryBe_1 = StoreBufferPlugin_hw_bypassQueryAddrIn[1 : 0];
  assign _zz__zz_StoreBufferPlugin_logic_loadQueryBe = ({3'd0,1'b1} <<< _zz_StoreBufferPlugin_logic_loadQueryBe_1);
  assign _zz__zz_StoreBufferPlugin_logic_loadQueryBe_2 = _zz__zz_StoreBufferPlugin_logic_loadQueryBe_3;
  assign _zz__zz_StoreBufferPlugin_logic_loadQueryBe_3 = ({3'd0,2'b11} <<< _zz__zz_StoreBufferPlugin_logic_loadQueryBe_4);
  assign _zz__zz_StoreBufferPlugin_logic_loadQueryBe_4 = ({1'd0,_zz_StoreBufferPlugin_logic_loadQueryBe_1[1 : 1]} <<< 1'd1);
  assign _zz__zz_StoreBufferPlugin_logic_loadQueryBe_5 = _zz__zz_StoreBufferPlugin_logic_loadQueryBe_6;
  assign _zz__zz_StoreBufferPlugin_logic_loadQueryBe_6 = ({3'd0,4'b1111} <<< 2'b00);
  assign _zz_FetchPipelinePlugin_logic_retryIdCounter_valueNext_1 = FetchPipelinePlugin_logic_retryIdCounter_willIncrement;
  assign _zz_FetchPipelinePlugin_logic_retryIdCounter_valueNext = {1'd0, _zz_FetchPipelinePlugin_logic_retryIdCounter_valueNext_1};
  assign _zz_FetchPipelinePlugin_logic_s2_logic_cmdPayload_transactionId = (s2_ICache_Access_FetchPipelinePlugin_logic_FetchPipeline_PC >>> 3'd4);
  assign _zz_219 = (s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC >>> 3'd4);
  assign _zz_218 = _zz_219[7:0];
  assign _zz__zz_io_push_payload_numValidInstructions = {1'd0, _zz_io_push_payload_numValidInstructions_2};
  assign _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag_1 = _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag[20 : 0];
  assign _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_1_tag = _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag[41 : 21];
  assign _zz__zz_ICachePlugin_logic_pipeline_f2_hitWayIdx = {ICachePlugin_logic_pipeline_f2_hit_ways_1,ICachePlugin_logic_pipeline_f2_hit_ways_0};
  assign _zz_ICachePlugin_logic_refill_refillCounter_valueNext_1 = ICachePlugin_logic_refill_refillCounter_willIncrement;
  assign _zz_ICachePlugin_logic_refill_refillCounter_valueNext = {1'd0, _zz_ICachePlugin_logic_refill_refillCounter_valueNext_1};
  assign _zz_io_uart_ar_bits_id = uartAxi_ar_payload_id;
  assign _zz_uartAxi_r_payload_id = io_uart_r_bits_id;
  assign _zz_io_uart_aw_bits_id = uartAxi_aw_payload_id;
  assign _zz_uartAxi_b_payload_id = io_uart_b_bits_id;
  assign _zz_io_leds_1 = (_zz_io_leds ? CommitPlugin_commitStatsReg_maxCommitPc : CommitPlugin_commitStatsReg_totalCommitted);
  assign _zz_ICachePlugin_logic_storage_tagLruRam_port = {ICachePlugin_logic_tag_write_logic_writeData_lru,{ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag,ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag}};
  assign _zz_ICachePlugin_logic_storage_dataRams_0_port = {ICachePlugin_logic_refill_lineBuffer_3,{ICachePlugin_logic_refill_lineBuffer_2,{ICachePlugin_logic_refill_lineBuffer_1,ICachePlugin_logic_refill_lineBuffer_0}}};
  assign _zz_ICachePlugin_logic_storage_dataRams_1_port = {ICachePlugin_logic_refill_lineBuffer_3,{ICachePlugin_logic_refill_lineBuffer_2,{ICachePlugin_logic_refill_lineBuffer_1,ICachePlugin_logic_refill_lineBuffer_0}}};
  assign _zz_BpuPipelinePlugin_logic_pht_port = BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_pc[11 : 2];
  assign _zz_BpuPipelinePlugin_logic_btb_port = BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_pc[9 : 2];
  assign _zz_BpuPipelinePlugin_logic_btb_port_1 = {BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_target,{BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_pc[31 : 10],1'b1}};
  assign _zz_CommitPlugin_logic_s0_committedThisCycle_comb_1 = CommitPlugin_logic_s0_commitAckMasks_0;
  assign _zz_CommitPlugin_logic_s0_recycledThisCycle_comb_1 = when_CommitPlugin_l265;
  assign _zz_DispatchPlugin_logic_destinationIqReady_4 = {_zz_DispatchPlugin_logic_destinationIqReady_2,_zz_DispatchPlugin_logic_destinationIqReady_1};
  assign _zz_DispatchPlugin_logic_dispatchOH = (s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_2_0_1);
  assign _zz_DispatchPlugin_logic_dispatchOH_1 = (s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_2_0_0);
  assign _zz_DispatchPlugin_logic_dispatchOH_2 = (s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_0_0_3);
  assign _zz_DispatchPlugin_logic_dispatchOH_3 = (s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_0_0_2);
  assign _zz_DispatchPlugin_logic_dispatchOH_4 = {(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_0_0_1),(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_0_0_0)};
  always @(posedge clk) begin
    if(ICachePlugin_logic_tag_write_logic_writeEnable) begin
      ICachePlugin_logic_storage_tagLruRam[ICachePlugin_logic_tag_write_logic_writeAddress] <= _zz_ICachePlugin_logic_storage_tagLruRam_port;
    end
  end

  always @(posedge clk) begin
    if(ICache_F1_Access_isFiring) begin
      ICachePlugin_logic_storage_tagLruRam_spinal_port1 <= ICachePlugin_logic_storage_tagLruRam[ICachePlugin_logic_pipeline_f1_f1_index];
    end
  end

  always @(posedge clk) begin
    if(ICache_F1_Access_isFiring) begin
      ICachePlugin_logic_storage_dataRams_0_spinal_port0 <= ICachePlugin_logic_storage_dataRams_0[ICachePlugin_logic_pipeline_f1_f1_index];
    end
  end

  always @(posedge clk) begin
    if(_zz_4) begin
      ICachePlugin_logic_storage_dataRams_0[_zz_ICachePlugin_logic_tag_write_logic_writeAddress] <= _zz_ICachePlugin_logic_storage_dataRams_0_port;
    end
  end

  always @(posedge clk) begin
    if(ICache_F1_Access_isFiring) begin
      ICachePlugin_logic_storage_dataRams_1_spinal_port0 <= ICachePlugin_logic_storage_dataRams_1[ICachePlugin_logic_pipeline_f1_f1_index];
    end
  end

  always @(posedge clk) begin
    if(_zz_3) begin
      ICachePlugin_logic_storage_dataRams_1[_zz_ICachePlugin_logic_tag_write_logic_writeAddress] <= _zz_ICachePlugin_logic_storage_dataRams_1_port;
    end
  end

  initial begin
    $readmemb("CoreNSCSCC.v_toplevel_BpuPipelinePlugin_logic_pht.bin",BpuPipelinePlugin_logic_pht);
  end
  always @(posedge clk) begin
    if(BpuPipelinePlugin_logic_s1_read_isFiring) begin
      BpuPipelinePlugin_logic_pht_spinal_port0 <= BpuPipelinePlugin_logic_pht[_zz_BpuPipelinePlugin_logic_phtReadData_s1];
    end
  end

  always @(posedge clk) begin
    if(BpuPipelinePlugin_logic_u1_read_isFiring) begin
      BpuPipelinePlugin_logic_pht_spinal_port1 <= BpuPipelinePlugin_logic_pht[_zz_BpuPipelinePlugin_logic_oldPhtState_u1];
    end
  end

  always @(posedge clk) begin
    if(_zz_2) begin
      BpuPipelinePlugin_logic_pht[_zz_BpuPipelinePlugin_logic_pht_port] <= BpuPipelinePlugin_logic_newPhtState;
    end
  end

  initial begin
    $readmemb("CoreNSCSCC.v_toplevel_BpuPipelinePlugin_logic_btb.bin",BpuPipelinePlugin_logic_btb);
  end
  always @(posedge clk) begin
    if(BpuPipelinePlugin_logic_s1_read_isFiring) begin
      BpuPipelinePlugin_logic_btb_spinal_port0 <= BpuPipelinePlugin_logic_btb[_zz_BpuPipelinePlugin_logic_btbReadData_s1_valid];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      BpuPipelinePlugin_logic_btb[_zz_BpuPipelinePlugin_logic_btb_port] <= _zz_BpuPipelinePlugin_logic_btb_port_1;
    end
  end

  IntAlu AluIntEU_AluIntEuPlugin_intAlu (
    .io_iqEntryIn_valid                          (s2_Execute_isFiring                                                  ), //i
    .io_iqEntryIn_payload_robPtr                 (_zz_io_iqEntryIn_payload_robPtr[3:0]                                 ), //i
    .io_iqEntryIn_payload_physDest_idx           (_zz_io_iqEntryIn_payload_physDest_idx[5:0]                           ), //i
    .io_iqEntryIn_payload_physDestIsFpr          (_zz_io_iqEntryIn_payload_physDestIsFpr                               ), //i
    .io_iqEntryIn_payload_writesToPhysReg        (_zz_io_iqEntryIn_payload_writesToPhysReg                             ), //i
    .io_iqEntryIn_payload_useSrc1                (_zz_io_iqEntryIn_payload_useSrc1                                     ), //i
    .io_iqEntryIn_payload_src1Data               (_zz_io_iqEntryIn_payload_src1Data[31:0]                              ), //i
    .io_iqEntryIn_payload_src1Tag                (_zz_io_iqEntryIn_payload_src1Tag[5:0]                                ), //i
    .io_iqEntryIn_payload_src1Ready              (_zz_io_iqEntryIn_payload_src1Ready                                   ), //i
    .io_iqEntryIn_payload_src1IsFpr              (_zz_io_iqEntryIn_payload_src1IsFpr                                   ), //i
    .io_iqEntryIn_payload_useSrc2                (_zz_io_iqEntryIn_payload_useSrc2                                     ), //i
    .io_iqEntryIn_payload_src2Data               (_zz_io_iqEntryIn_payload_src2Data_1[31:0]                            ), //i
    .io_iqEntryIn_payload_src2Tag                (_zz_io_iqEntryIn_payload_src2Tag[5:0]                                ), //i
    .io_iqEntryIn_payload_src2Ready              (_zz_io_iqEntryIn_payload_src2Ready                                   ), //i
    .io_iqEntryIn_payload_src2IsFpr              (_zz_io_iqEntryIn_payload_src2IsFpr                                   ), //i
    .io_iqEntryIn_payload_aluCtrl_valid          (_zz_io_iqEntryIn_payload_aluCtrl_valid                               ), //i
    .io_iqEntryIn_payload_aluCtrl_isSub          (_zz_io_iqEntryIn_payload_aluCtrl_isSub                               ), //i
    .io_iqEntryIn_payload_aluCtrl_isAdd          (_zz_io_iqEntryIn_payload_aluCtrl_isAdd                               ), //i
    .io_iqEntryIn_payload_aluCtrl_isSigned       (_zz_io_iqEntryIn_payload_aluCtrl_isSigned                            ), //i
    .io_iqEntryIn_payload_aluCtrl_logicOp        (_zz_io_iqEntryIn_payload_aluCtrl_logicOp[1:0]                        ), //i
    .io_iqEntryIn_payload_shiftCtrl_valid        (_zz_io_iqEntryIn_payload_shiftCtrl_valid                             ), //i
    .io_iqEntryIn_payload_shiftCtrl_isRight      (_zz_io_iqEntryIn_payload_shiftCtrl_isRight                           ), //i
    .io_iqEntryIn_payload_shiftCtrl_isArithmetic (_zz_io_iqEntryIn_payload_shiftCtrl_isArithmetic                      ), //i
    .io_iqEntryIn_payload_shiftCtrl_isRotate     (_zz_io_iqEntryIn_payload_shiftCtrl_isRotate                          ), //i
    .io_iqEntryIn_payload_shiftCtrl_isDoubleWord (_zz_io_iqEntryIn_payload_shiftCtrl_isDoubleWord                      ), //i
    .io_iqEntryIn_payload_imm                    (_zz_io_iqEntryIn_payload_imm[31:0]                                   ), //i
    .io_iqEntryIn_payload_immUsage               (_zz_io_iqEntryIn_payload_immUsage[2:0]                               ), //i
    .io_resultOut_valid                          (AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_valid                    ), //o
    .io_resultOut_payload_data                   (AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_data[31:0]       ), //o
    .io_resultOut_payload_physDest_idx           (AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_physDest_idx[5:0]), //o
    .io_resultOut_payload_writesToPhysReg        (AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_writesToPhysReg  ), //o
    .io_resultOut_payload_robPtr                 (AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_robPtr[3:0]      ), //o
    .io_resultOut_payload_hasException           (AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_hasException     ), //o
    .io_resultOut_payload_exceptionCode          (AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_exceptionCode    )  //o
  );
  SRAMController CoreMemSysPlugin_hw_baseramCtrl (
    .io_axi_aw_valid         (axi4WriteOnlyArbiter_3_io_output_aw_valid                  ), //i
    .io_axi_aw_ready         (CoreMemSysPlugin_hw_baseramCtrl_io_axi_aw_ready            ), //o
    .io_axi_aw_payload_addr  (axi4WriteOnlyArbiter_3_io_output_aw_payload_addr[31:0]     ), //i
    .io_axi_aw_payload_id    (axi4WriteOnlyArbiter_3_io_output_aw_payload_id[6:0]        ), //i
    .io_axi_aw_payload_len   (axi4WriteOnlyArbiter_3_io_output_aw_payload_len[7:0]       ), //i
    .io_axi_aw_payload_size  (axi4WriteOnlyArbiter_3_io_output_aw_payload_size[2:0]      ), //i
    .io_axi_aw_payload_burst (axi4WriteOnlyArbiter_3_io_output_aw_payload_burst[1:0]     ), //i
    .io_axi_w_valid          (axi4WriteOnlyArbiter_3_io_output_w_valid                   ), //i
    .io_axi_w_ready          (CoreMemSysPlugin_hw_baseramCtrl_io_axi_w_ready             ), //o
    .io_axi_w_payload_data   (axi4WriteOnlyArbiter_3_io_output_w_payload_data[31:0]      ), //i
    .io_axi_w_payload_strb   (axi4WriteOnlyArbiter_3_io_output_w_payload_strb[3:0]       ), //i
    .io_axi_w_payload_last   (axi4WriteOnlyArbiter_3_io_output_w_payload_last            ), //i
    .io_axi_b_valid          (CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_valid             ), //o
    .io_axi_b_ready          (axi4WriteOnlyArbiter_3_io_output_b_ready                   ), //i
    .io_axi_b_payload_id     (CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_payload_id[6:0]   ), //o
    .io_axi_b_payload_resp   (CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_payload_resp[1:0] ), //o
    .io_axi_ar_valid         (axi4ReadOnlyArbiter_3_io_output_ar_valid                   ), //i
    .io_axi_ar_ready         (CoreMemSysPlugin_hw_baseramCtrl_io_axi_ar_ready            ), //o
    .io_axi_ar_payload_addr  (axi4ReadOnlyArbiter_3_io_output_ar_payload_addr[31:0]      ), //i
    .io_axi_ar_payload_id    (axi4ReadOnlyArbiter_3_io_output_ar_payload_id[6:0]         ), //i
    .io_axi_ar_payload_len   (axi4ReadOnlyArbiter_3_io_output_ar_payload_len[7:0]        ), //i
    .io_axi_ar_payload_size  (axi4ReadOnlyArbiter_3_io_output_ar_payload_size[2:0]       ), //i
    .io_axi_ar_payload_burst (axi4ReadOnlyArbiter_3_io_output_ar_payload_burst[1:0]      ), //i
    .io_axi_r_valid          (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_valid             ), //o
    .io_axi_r_ready          (axi4ReadOnlyArbiter_3_io_output_r_ready                    ), //i
    .io_axi_r_payload_data   (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_data[31:0]), //o
    .io_axi_r_payload_id     (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_id[6:0]   ), //o
    .io_axi_r_payload_resp   (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_resp[1:0] ), //o
    .io_axi_r_payload_last   (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_last      ), //o
    .io_ram_data_read        (io_isram_dout[31:0]                                        ), //i
    .io_ram_data_write       (CoreMemSysPlugin_hw_baseramCtrl_io_ram_data_write[31:0]    ), //o
    .io_ram_data_writeEnable (CoreMemSysPlugin_hw_baseramCtrl_io_ram_data_writeEnable    ), //o
    .io_ram_addr             (CoreMemSysPlugin_hw_baseramCtrl_io_ram_addr[19:0]          ), //o
    .io_ram_be_n             (CoreMemSysPlugin_hw_baseramCtrl_io_ram_be_n[3:0]           ), //o
    .io_ram_ce_n             (CoreMemSysPlugin_hw_baseramCtrl_io_ram_ce_n                ), //o
    .io_ram_oe_n             (CoreMemSysPlugin_hw_baseramCtrl_io_ram_oe_n                ), //o
    .io_ram_we_n             (CoreMemSysPlugin_hw_baseramCtrl_io_ram_we_n                ), //o
    .clk                     (clk                                                        ), //i
    .reset                   (reset                                                      )  //i
  );
  SRAMController_1 CoreMemSysPlugin_hw_extramCtrl (
    .io_axi_aw_valid         (axi4WriteOnlyArbiter_4_io_output_aw_valid                 ), //i
    .io_axi_aw_ready         (CoreMemSysPlugin_hw_extramCtrl_io_axi_aw_ready            ), //o
    .io_axi_aw_payload_addr  (axi4WriteOnlyArbiter_4_io_output_aw_payload_addr[31:0]    ), //i
    .io_axi_aw_payload_id    (axi4WriteOnlyArbiter_4_io_output_aw_payload_id[6:0]       ), //i
    .io_axi_aw_payload_len   (axi4WriteOnlyArbiter_4_io_output_aw_payload_len[7:0]      ), //i
    .io_axi_aw_payload_size  (axi4WriteOnlyArbiter_4_io_output_aw_payload_size[2:0]     ), //i
    .io_axi_aw_payload_burst (axi4WriteOnlyArbiter_4_io_output_aw_payload_burst[1:0]    ), //i
    .io_axi_w_valid          (axi4WriteOnlyArbiter_4_io_output_w_valid                  ), //i
    .io_axi_w_ready          (CoreMemSysPlugin_hw_extramCtrl_io_axi_w_ready             ), //o
    .io_axi_w_payload_data   (axi4WriteOnlyArbiter_4_io_output_w_payload_data[31:0]     ), //i
    .io_axi_w_payload_strb   (axi4WriteOnlyArbiter_4_io_output_w_payload_strb[3:0]      ), //i
    .io_axi_w_payload_last   (axi4WriteOnlyArbiter_4_io_output_w_payload_last           ), //i
    .io_axi_b_valid          (CoreMemSysPlugin_hw_extramCtrl_io_axi_b_valid             ), //o
    .io_axi_b_ready          (axi4WriteOnlyArbiter_4_io_output_b_ready                  ), //i
    .io_axi_b_payload_id     (CoreMemSysPlugin_hw_extramCtrl_io_axi_b_payload_id[6:0]   ), //o
    .io_axi_b_payload_resp   (CoreMemSysPlugin_hw_extramCtrl_io_axi_b_payload_resp[1:0] ), //o
    .io_axi_ar_valid         (axi4ReadOnlyArbiter_4_io_output_ar_valid                  ), //i
    .io_axi_ar_ready         (CoreMemSysPlugin_hw_extramCtrl_io_axi_ar_ready            ), //o
    .io_axi_ar_payload_addr  (axi4ReadOnlyArbiter_4_io_output_ar_payload_addr[31:0]     ), //i
    .io_axi_ar_payload_id    (axi4ReadOnlyArbiter_4_io_output_ar_payload_id[6:0]        ), //i
    .io_axi_ar_payload_len   (axi4ReadOnlyArbiter_4_io_output_ar_payload_len[7:0]       ), //i
    .io_axi_ar_payload_size  (axi4ReadOnlyArbiter_4_io_output_ar_payload_size[2:0]      ), //i
    .io_axi_ar_payload_burst (axi4ReadOnlyArbiter_4_io_output_ar_payload_burst[1:0]     ), //i
    .io_axi_r_valid          (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_valid             ), //o
    .io_axi_r_ready          (axi4ReadOnlyArbiter_4_io_output_r_ready                   ), //i
    .io_axi_r_payload_data   (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_data[31:0]), //o
    .io_axi_r_payload_id     (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_id[6:0]   ), //o
    .io_axi_r_payload_resp   (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_resp[1:0] ), //o
    .io_axi_r_payload_last   (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_last      ), //o
    .io_ram_data_read        (io_dsram_dout[31:0]                                       ), //i
    .io_ram_data_write       (CoreMemSysPlugin_hw_extramCtrl_io_ram_data_write[31:0]    ), //o
    .io_ram_data_writeEnable (CoreMemSysPlugin_hw_extramCtrl_io_ram_data_writeEnable    ), //o
    .io_ram_addr             (CoreMemSysPlugin_hw_extramCtrl_io_ram_addr[19:0]          ), //o
    .io_ram_be_n             (CoreMemSysPlugin_hw_extramCtrl_io_ram_be_n[3:0]           ), //o
    .io_ram_ce_n             (CoreMemSysPlugin_hw_extramCtrl_io_ram_ce_n                ), //o
    .io_ram_oe_n             (CoreMemSysPlugin_hw_extramCtrl_io_ram_oe_n                ), //o
    .io_ram_we_n             (CoreMemSysPlugin_hw_extramCtrl_io_ram_we_n                ), //o
    .clk                     (clk                                                       ), //i
    .reset                   (reset                                                     )  //i
  );
  DataCache DataCachePlugin_setup_cache (
    .io_load_cmd_valid                         (DataCachePlugin_logic_load_hit                                             ), //i
    .io_load_cmd_ready                         (DataCachePlugin_setup_cache_io_load_cmd_ready                              ), //o
    .io_load_cmd_payload_virtual               (LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_virtual[31:0]                ), //i
    .io_load_cmd_payload_size                  (LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size[1:0]                    ), //i
    .io_load_cmd_payload_redoOnDataHazard      (LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_redoOnDataHazard             ), //i
    .io_load_cmd_payload_transactionId         (LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_transactionId[2:0]           ), //i
    .io_load_cmd_payload_id                    (LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_id[2:0]                      ), //i
    .io_load_translated_physical               (LoadQueuePlugin_hw_dCacheLoadPort_translated_physical[31:0]                ), //i
    .io_load_translated_abord                  (LoadQueuePlugin_hw_dCacheLoadPort_translated_abord                         ), //i
    .io_load_cancels                           (LoadQueuePlugin_hw_dCacheLoadPort_cancels[2:0]                             ), //i
    .io_load_rsp_valid                         (DataCachePlugin_setup_cache_io_load_rsp_valid                              ), //o
    .io_load_rsp_payload_data                  (DataCachePlugin_setup_cache_io_load_rsp_payload_data[31:0]                 ), //o
    .io_load_rsp_payload_fault                 (DataCachePlugin_setup_cache_io_load_rsp_payload_fault                      ), //o
    .io_load_rsp_payload_redo                  (DataCachePlugin_setup_cache_io_load_rsp_payload_redo                       ), //o
    .io_load_rsp_payload_refillSlot            (DataCachePlugin_setup_cache_io_load_rsp_payload_refillSlot[7:0]            ), //o
    .io_load_rsp_payload_refillSlotAny         (DataCachePlugin_setup_cache_io_load_rsp_payload_refillSlotAny              ), //o
    .io_load_rsp_payload_id                    (DataCachePlugin_setup_cache_io_load_rsp_payload_id[2:0]                    ), //o
    .io_store_cmd_valid                        (StoreBufferPlugin_hw_dCacheStorePort_cmd_valid                             ), //i
    .io_store_cmd_ready                        (DataCachePlugin_setup_cache_io_store_cmd_ready                             ), //o
    .io_store_cmd_payload_address              (StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_address[31:0]             ), //i
    .io_store_cmd_payload_data                 (StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_data[31:0]                ), //i
    .io_store_cmd_payload_mask                 (StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_mask[3:0]                 ), //i
    .io_store_cmd_payload_io                   (StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_io                        ), //i
    .io_store_cmd_payload_flush                (StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flush                     ), //i
    .io_store_cmd_payload_flushFree            (StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flushFree                 ), //i
    .io_store_cmd_payload_prefetch             (StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_prefetch                  ), //i
    .io_store_cmd_payload_id                   (StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_id[2:0]                   ), //i
    .io_store_rsp_valid                        (DataCachePlugin_setup_cache_io_store_rsp_valid                             ), //o
    .io_store_rsp_payload_fault                (DataCachePlugin_setup_cache_io_store_rsp_payload_fault                     ), //o
    .io_store_rsp_payload_redo                 (DataCachePlugin_setup_cache_io_store_rsp_payload_redo                      ), //o
    .io_store_rsp_payload_refillSlot           (DataCachePlugin_setup_cache_io_store_rsp_payload_refillSlot[7:0]           ), //o
    .io_store_rsp_payload_refillSlotAny        (DataCachePlugin_setup_cache_io_store_rsp_payload_refillSlotAny             ), //o
    .io_store_rsp_payload_flush                (DataCachePlugin_setup_cache_io_store_rsp_payload_flush                     ), //o
    .io_store_rsp_payload_prefetch             (DataCachePlugin_setup_cache_io_store_rsp_payload_prefetch                  ), //o
    .io_store_rsp_payload_address              (DataCachePlugin_setup_cache_io_store_rsp_payload_address[31:0]             ), //o
    .io_store_rsp_payload_io                   (DataCachePlugin_setup_cache_io_store_rsp_payload_io                        ), //o
    .io_store_rsp_payload_id                   (DataCachePlugin_setup_cache_io_store_rsp_payload_id[2:0]                   ), //o
    .io_mem_read_cmd_valid                     (DataCachePlugin_setup_cache_io_mem_read_cmd_valid                          ), //o
    .io_mem_read_cmd_ready                     (DataCachePlugin_setup_cache_io_mem_read_cmd_ready                          ), //i
    .io_mem_read_cmd_payload_id                (DataCachePlugin_setup_cache_io_mem_read_cmd_payload_id[2:0]                ), //o
    .io_mem_read_cmd_payload_address           (DataCachePlugin_setup_cache_io_mem_read_cmd_payload_address[31:0]          ), //o
    .io_mem_read_rsp_valid                     (io_mem_toAxi4_rRspStaged_valid                                             ), //i
    .io_mem_read_rsp_ready                     (DataCachePlugin_setup_cache_io_mem_read_rsp_ready                          ), //o
    .io_mem_read_rsp_payload_id                (io_mem_toAxi4_rRspStaged_payload_id[2:0]                                   ), //i
    .io_mem_read_rsp_payload_data              (io_mem_toAxi4_rRspStaged_payload_data[31:0]                                ), //i
    .io_mem_read_rsp_payload_error             (DataCachePlugin_setup_cache_io_mem_read_rsp_payload_error                  ), //i
    .io_mem_write_cmd_valid                    (DataCachePlugin_setup_cache_io_mem_write_cmd_valid                         ), //o
    .io_mem_write_cmd_ready                    (DataCachePlugin_setup_cache_io_mem_write_cmd_ready                         ), //i
    .io_mem_write_cmd_payload_last             (DataCachePlugin_setup_cache_io_mem_write_cmd_payload_last                  ), //o
    .io_mem_write_cmd_payload_fragment_address (DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_address[31:0]), //o
    .io_mem_write_cmd_payload_fragment_data    (DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_data[31:0]   ), //o
    .io_mem_write_cmd_payload_fragment_id      (DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_id[2:0]      ), //o
    .io_mem_write_rsp_valid                    (io_mem_toAxi4_bRspStaged_valid                                             ), //i
    .io_mem_write_rsp_payload_error            (DataCachePlugin_setup_cache_io_mem_write_rsp_payload_error                 ), //i
    .io_mem_write_rsp_payload_id               (io_mem_toAxi4_bRspStaged_payload_id[2:0]                                   ), //i
    .io_refillCompletions                      (DataCachePlugin_setup_cache_io_refillCompletions[7:0]                      ), //o
    .io_refillEvent                            (DataCachePlugin_setup_cache_io_refillEvent                                 ), //o
    .io_writebackEvent                         (DataCachePlugin_setup_cache_io_writebackEvent                              ), //o
    .io_writebackBusy                          (DataCachePlugin_setup_cache_io_writebackBusy                               ), //o
    .clk                                       (clk                                                                        ), //i
    .reset                                     (reset                                                                      )  //i
  );
  OneShot oneShot_13 (
    .io_triggerIn (oneShot_13_io_triggerIn), //i
    .io_pulseOut  (oneShot_13_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  StreamFifo_11 FetchPipelinePlugin_setup_fetchOutput (
    .io_push_valid                              (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_valid                             ), //i
    .io_push_ready                              (FetchPipelinePlugin_setup_fetchOutput_io_push_ready                                   ), //o
    .io_push_payload_pc                         (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_pc[31:0]                  ), //i
    .io_push_payload_instruction                (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_instruction[31:0]         ), //i
    .io_push_payload_predecode_isBranch         (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isBranch        ), //i
    .io_push_payload_predecode_isJump           (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isJump          ), //i
    .io_push_payload_predecode_isDirectJump     (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isDirectJump    ), //i
    .io_push_payload_predecode_jumpOffset       (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_jumpOffset[31:0]), //i
    .io_push_payload_predecode_isIdle           (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isIdle          ), //i
    .io_push_payload_bpuPrediction_isTaken      (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_isTaken     ), //i
    .io_push_payload_bpuPrediction_target       (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_target[31:0]), //i
    .io_push_payload_bpuPrediction_wasPredicted (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_wasPredicted), //i
    .io_pop_valid                               (FetchPipelinePlugin_setup_fetchOutput_io_pop_valid                                    ), //o
    .io_pop_ready                               (s0_Decode_ready                                                                       ), //i
    .io_pop_payload_pc                          (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_pc[31:0]                         ), //o
    .io_pop_payload_instruction                 (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_instruction[31:0]                ), //o
    .io_pop_payload_predecode_isBranch          (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_isBranch               ), //o
    .io_pop_payload_predecode_isJump            (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_isJump                 ), //o
    .io_pop_payload_predecode_isDirectJump      (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_isDirectJump           ), //o
    .io_pop_payload_predecode_jumpOffset        (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_jumpOffset[31:0]       ), //o
    .io_pop_payload_predecode_isIdle            (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_predecode_isIdle                 ), //o
    .io_pop_payload_bpuPrediction_isTaken       (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_isTaken            ), //o
    .io_pop_payload_bpuPrediction_target        (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_target[31:0]       ), //o
    .io_pop_payload_bpuPrediction_wasPredicted  (FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_wasPredicted       ), //o
    .io_flush                                   (FetchPipelinePlugin_logic_hardRedirect_valid                                          ), //i
    .io_occupancy                               (FetchPipelinePlugin_setup_fetchOutput_io_occupancy[2:0]                               ), //o
    .io_availability                            (FetchPipelinePlugin_setup_fetchOutput_io_availability[2:0]                            ), //o
    .clk                                        (clk                                                                                   ), //i
    .reset                                      (reset                                                                                 )  //i
  );
  ReorderBuffer ROBPlugin_robComponent (
    .io_allocate_0_valid                                                 (ROBPlugin_robComponent_io_allocate_0_valid                                                ), //i
    .io_allocate_0_uopIn_decoded_pc                                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_pc[31:0]                          ), //i
    .io_allocate_0_uopIn_decoded_isValid                                 (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isValid                           ), //i
    .io_allocate_0_uopIn_decoded_uopCode                                 (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode[4:0]                      ), //i
    .io_allocate_0_uopIn_decoded_exeUnit                                 (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit[3:0]                      ), //i
    .io_allocate_0_uopIn_decoded_isa                                     (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa[1:0]                          ), //i
    .io_allocate_0_uopIn_decoded_archDest_idx                            (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_idx[4:0]                 ), //i
    .io_allocate_0_uopIn_decoded_archDest_rtype                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype[1:0]               ), //i
    .io_allocate_0_uopIn_decoded_writeArchDestEn                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_writeArchDestEn                   ), //i
    .io_allocate_0_uopIn_decoded_archSrc1_idx                            (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_idx[4:0]                 ), //i
    .io_allocate_0_uopIn_decoded_archSrc1_rtype                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype[1:0]               ), //i
    .io_allocate_0_uopIn_decoded_useArchSrc1                             (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_useArchSrc1                       ), //i
    .io_allocate_0_uopIn_decoded_archSrc2_idx                            (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_idx[4:0]                 ), //i
    .io_allocate_0_uopIn_decoded_archSrc2_rtype                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype[1:0]               ), //i
    .io_allocate_0_uopIn_decoded_useArchSrc2                             (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_useArchSrc2                       ), //i
    .io_allocate_0_uopIn_decoded_usePcForAddr                            (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_usePcForAddr                      ), //i
    .io_allocate_0_uopIn_decoded_imm                                     (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_imm[31:0]                         ), //i
    .io_allocate_0_uopIn_decoded_immUsage                                (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage[2:0]                     ), //i
    .io_allocate_0_uopIn_decoded_aluCtrl_valid                           (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_valid                     ), //i
    .io_allocate_0_uopIn_decoded_aluCtrl_isSub                           (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isSub                     ), //i
    .io_allocate_0_uopIn_decoded_aluCtrl_isAdd                           (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isAdd                     ), //i
    .io_allocate_0_uopIn_decoded_aluCtrl_isSigned                        (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isSigned                  ), //i
    .io_allocate_0_uopIn_decoded_aluCtrl_logicOp                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp[1:0]              ), //i
    .io_allocate_0_uopIn_decoded_shiftCtrl_valid                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_valid                   ), //i
    .io_allocate_0_uopIn_decoded_shiftCtrl_isRight                       (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isRight                 ), //i
    .io_allocate_0_uopIn_decoded_shiftCtrl_isArithmetic                  (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isArithmetic            ), //i
    .io_allocate_0_uopIn_decoded_shiftCtrl_isRotate                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isRotate                ), //i
    .io_allocate_0_uopIn_decoded_shiftCtrl_isDoubleWord                  (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isDoubleWord            ), //i
    .io_allocate_0_uopIn_decoded_mulDivCtrl_valid                        (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_valid                  ), //i
    .io_allocate_0_uopIn_decoded_mulDivCtrl_isDiv                        (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isDiv                  ), //i
    .io_allocate_0_uopIn_decoded_mulDivCtrl_isSigned                     (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isSigned               ), //i
    .io_allocate_0_uopIn_decoded_mulDivCtrl_isWordOp                     (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isWordOp               ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_size                            (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size[1:0]                 ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_isSignedLoad                    (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isSignedLoad              ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_isStore                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isStore                   ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_isLoadLinked                    (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isLoadLinked              ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_isStoreCond                     (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isStoreCond               ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_atomicOp                        (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_atomicOp[4:0]             ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_isFence                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isFence                   ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_fenceMode                       (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_fenceMode[7:0]            ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_isCacheOp                       (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isCacheOp                 ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_cacheOpType                     (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_cacheOpType[4:0]          ), //i
    .io_allocate_0_uopIn_decoded_memCtrl_isPrefetch                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isPrefetch                ), //i
    .io_allocate_0_uopIn_decoded_branchCtrl_condition                    (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition[4:0]         ), //i
    .io_allocate_0_uopIn_decoded_branchCtrl_isJump                       (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isJump                 ), //i
    .io_allocate_0_uopIn_decoded_branchCtrl_isLink                       (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isLink                 ), //i
    .io_allocate_0_uopIn_decoded_branchCtrl_linkReg_idx                  (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_idx[4:0]       ), //i
    .io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype                (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype[1:0]     ), //i
    .io_allocate_0_uopIn_decoded_branchCtrl_isIndirect                   (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isIndirect             ), //i
    .io_allocate_0_uopIn_decoded_branchCtrl_laCfIdx                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_laCfIdx[2:0]           ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_opType                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_opType[3:0]               ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1[1:0]           ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2[1:0]           ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest[1:0]           ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_roundingMode                    (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_roundingMode[2:0]         ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_isIntegerDest                   (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_isIntegerDest             ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_isSignedCvt                     (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_isSignedCvt               ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_fmaNegSrc1                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1                ), //i
    .io_allocate_0_uopIn_decoded_fpuCtrl_fcmpCond                        (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fcmpCond[4:0]             ), //i
    .io_allocate_0_uopIn_decoded_csrCtrl_csrAddr                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_csrAddr[13:0]             ), //i
    .io_allocate_0_uopIn_decoded_csrCtrl_isWrite                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isWrite                   ), //i
    .io_allocate_0_uopIn_decoded_csrCtrl_isRead                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isRead                    ), //i
    .io_allocate_0_uopIn_decoded_csrCtrl_isExchange                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isExchange                ), //i
    .io_allocate_0_uopIn_decoded_csrCtrl_useUimmAsSrc                    (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_useUimmAsSrc              ), //i
    .io_allocate_0_uopIn_decoded_sysCtrl_sysCode                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_sysCode[19:0]             ), //i
    .io_allocate_0_uopIn_decoded_sysCtrl_isExceptionReturn               (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_isExceptionReturn         ), //i
    .io_allocate_0_uopIn_decoded_sysCtrl_isTlbOp                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_isTlbOp                   ), //i
    .io_allocate_0_uopIn_decoded_sysCtrl_tlbOpType                       (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_tlbOpType[3:0]            ), //i
    .io_allocate_0_uopIn_decoded_decodeExceptionCode                     (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode[1:0]          ), //i
    .io_allocate_0_uopIn_decoded_hasDecodeException                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_hasDecodeException                ), //i
    .io_allocate_0_uopIn_decoded_isMicrocode                             (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isMicrocode                       ), //i
    .io_allocate_0_uopIn_decoded_microcodeEntry                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_microcodeEntry[7:0]               ), //i
    .io_allocate_0_uopIn_decoded_isSerializing                           (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isSerializing                     ), //i
    .io_allocate_0_uopIn_decoded_isBranchOrJump                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isBranchOrJump                    ), //i
    .io_allocate_0_uopIn_decoded_branchPrediction_isTaken                (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_isTaken          ), //i
    .io_allocate_0_uopIn_decoded_branchPrediction_target                 (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_target[31:0]     ), //i
    .io_allocate_0_uopIn_decoded_branchPrediction_wasPredicted           (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_wasPredicted     ), //i
    .io_allocate_0_uopIn_rename_physSrc1_idx                             (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc1_idx[5:0]                  ), //i
    .io_allocate_0_uopIn_rename_physSrc1IsFpr                            (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc1IsFpr                      ), //i
    .io_allocate_0_uopIn_rename_physSrc2_idx                             (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc2_idx[5:0]                  ), //i
    .io_allocate_0_uopIn_rename_physSrc2IsFpr                            (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc2IsFpr                      ), //i
    .io_allocate_0_uopIn_rename_physDest_idx                             (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physDest_idx[5:0]                  ), //i
    .io_allocate_0_uopIn_rename_physDestIsFpr                            (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physDestIsFpr                      ), //i
    .io_allocate_0_uopIn_rename_oldPhysDest_idx                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_oldPhysDest_idx[5:0]               ), //i
    .io_allocate_0_uopIn_rename_oldPhysDestIsFpr                         (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_oldPhysDestIsFpr                   ), //i
    .io_allocate_0_uopIn_rename_allocatesPhysDest                        (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_allocatesPhysDest                  ), //i
    .io_allocate_0_uopIn_rename_writesToPhysReg                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_writesToPhysReg                    ), //i
    .io_allocate_0_uopIn_robPtr                                          (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_robPtr[3:0]                               ), //i
    .io_allocate_0_uopIn_uniqueId                                        (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_uniqueId[15:0]                            ), //i
    .io_allocate_0_uopIn_dispatched                                      (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_dispatched                                ), //i
    .io_allocate_0_uopIn_executed                                        (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_executed                                  ), //i
    .io_allocate_0_uopIn_hasException                                    (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_hasException                              ), //i
    .io_allocate_0_uopIn_exceptionCode                                   (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_exceptionCode[7:0]                        ), //i
    .io_allocate_0_pcIn                                                  (s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_pc[31:0]                          ), //i
    .io_allocate_0_robPtr                                                (ROBPlugin_robComponent_io_allocate_0_robPtr[3:0]                                          ), //o
    .io_allocate_0_ready                                                 (ROBPlugin_robComponent_io_allocate_0_ready                                                ), //o
    .io_canAllocate_0                                                    (ROBPlugin_robComponent_io_canAllocate_0                                                   ), //o
    .io_writeback_0_fire                                                 (AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes                                     ), //i
    .io_writeback_0_robPtr                                               (AluIntEU_AluIntEuPlugin_euResult_uop_robPtr[3:0]                                          ), //i
    .io_writeback_0_isTaken                                              (AluIntEU_AluIntEuPlugin_euResult_isTaken                                                  ), //i
    .io_writeback_0_isMispredictedBranch                                 (AluIntEU_AluIntEuPlugin_euResult_isMispredictedBranch                                     ), //i
    .io_writeback_0_result                                               (AluIntEU_AluIntEuPlugin_euResult_data[31:0]                                               ), //i
    .io_writeback_0_exceptionOccurred                                    (AluIntEU_AluIntEuPlugin_euResult_hasException                                             ), //i
    .io_writeback_0_exceptionCodeIn                                      (AluIntEU_AluIntEuPlugin_euResult_exceptionCode[7:0]                                       ), //i
    .io_writeback_1_fire                                                 (MulEU_MulEuPlugin_logicPhase_executionCompletes                                           ), //i
    .io_writeback_1_robPtr                                               (MulEU_MulEuPlugin_euResult_uop_robPtr[3:0]                                                ), //i
    .io_writeback_1_isTaken                                              (MulEU_MulEuPlugin_euResult_isTaken                                                        ), //i
    .io_writeback_1_isMispredictedBranch                                 (MulEU_MulEuPlugin_euResult_isMispredictedBranch                                           ), //i
    .io_writeback_1_result                                               (MulEU_MulEuPlugin_euResult_data[31:0]                                                     ), //i
    .io_writeback_1_exceptionOccurred                                    (MulEU_MulEuPlugin_euResult_hasException                                                   ), //i
    .io_writeback_1_exceptionCodeIn                                      (MulEU_MulEuPlugin_euResult_exceptionCode[7:0]                                             ), //i
    .io_writeback_2_fire                                                 (BranchEU_BranchEuPlugin_logicPhase_executionCompletes                                     ), //i
    .io_writeback_2_robPtr                                               (BranchEU_BranchEuPlugin_euResult_uop_robPtr[3:0]                                          ), //i
    .io_writeback_2_isTaken                                              (BranchEU_BranchEuPlugin_euResult_isTaken                                                  ), //i
    .io_writeback_2_isMispredictedBranch                                 (BranchEU_BranchEuPlugin_euResult_isMispredictedBranch                                     ), //i
    .io_writeback_2_result                                               (BranchEU_BranchEuPlugin_euResult_data[31:0]                                               ), //i
    .io_writeback_2_exceptionOccurred                                    (BranchEU_BranchEuPlugin_euResult_hasException                                             ), //i
    .io_writeback_2_exceptionCodeIn                                      (BranchEU_BranchEuPlugin_euResult_exceptionCode[7:0]                                       ), //i
    .io_writeback_3_fire                                                 (LsuEU_LsuEuPlugin_logicPhase_executionCompletes                                           ), //i
    .io_writeback_3_robPtr                                               (LsuEU_LsuEuPlugin_euResult_uop_robPtr[3:0]                                                ), //i
    .io_writeback_3_isTaken                                              (LsuEU_LsuEuPlugin_euResult_isTaken                                                        ), //i
    .io_writeback_3_isMispredictedBranch                                 (LsuEU_LsuEuPlugin_euResult_isMispredictedBranch                                           ), //i
    .io_writeback_3_result                                               (LsuEU_LsuEuPlugin_euResult_data[31:0]                                                     ), //i
    .io_writeback_3_exceptionOccurred                                    (LsuEU_LsuEuPlugin_euResult_hasException                                                   ), //i
    .io_writeback_3_exceptionCodeIn                                      (LsuEU_LsuEuPlugin_euResult_exceptionCode[7:0]                                             ), //i
    .io_writeback_4_fire                                                 (ROBPlugin_robComponent_io_writeback_4_fire                                                ), //i
    .io_writeback_4_robPtr                                               (ROBPlugin_robComponent_io_writeback_4_robPtr[3:0]                                         ), //i
    .io_writeback_4_isTaken                                              (1'bx                                                                                      ), //i
    .io_writeback_4_isMispredictedBranch                                 (1'bx                                                                                      ), //i
    .io_writeback_4_result                                               (ROBPlugin_robComponent_io_writeback_4_result[31:0]                                        ), //i
    .io_writeback_4_exceptionOccurred                                    (ROBPlugin_robComponent_io_writeback_4_exceptionOccurred                                   ), //i
    .io_writeback_4_exceptionCodeIn                                      (ROBPlugin_robComponent_io_writeback_4_exceptionCodeIn[7:0]                                ), //i
    .io_commit_0_valid                                                   (ROBPlugin_robComponent_io_commit_0_valid                                                  ), //o
    .io_commit_0_canCommit                                               (ROBPlugin_robComponent_io_commit_0_canCommit                                              ), //o
    .io_commit_0_entry_payload_uop_decoded_pc                            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_pc[31:0]                     ), //o
    .io_commit_0_entry_payload_uop_decoded_isValid                       (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isValid                      ), //o
    .io_commit_0_entry_payload_uop_decoded_uopCode                       (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_uopCode[4:0]                 ), //o
    .io_commit_0_entry_payload_uop_decoded_exeUnit                       (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_exeUnit[3:0]                 ), //o
    .io_commit_0_entry_payload_uop_decoded_isa                           (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isa[1:0]                     ), //o
    .io_commit_0_entry_payload_uop_decoded_archDest_idx                  (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archDest_idx[4:0]            ), //o
    .io_commit_0_entry_payload_uop_decoded_archDest_rtype                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archDest_rtype[1:0]          ), //o
    .io_commit_0_entry_payload_uop_decoded_writeArchDestEn               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_writeArchDestEn              ), //o
    .io_commit_0_entry_payload_uop_decoded_archSrc1_idx                  (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archSrc1_idx[4:0]            ), //o
    .io_commit_0_entry_payload_uop_decoded_archSrc1_rtype                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype[1:0]          ), //o
    .io_commit_0_entry_payload_uop_decoded_useArchSrc1                   (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_useArchSrc1                  ), //o
    .io_commit_0_entry_payload_uop_decoded_archSrc2_idx                  (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archSrc2_idx[4:0]            ), //o
    .io_commit_0_entry_payload_uop_decoded_archSrc2_rtype                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype[1:0]          ), //o
    .io_commit_0_entry_payload_uop_decoded_useArchSrc2                   (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_useArchSrc2                  ), //o
    .io_commit_0_entry_payload_uop_decoded_usePcForAddr                  (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_usePcForAddr                 ), //o
    .io_commit_0_entry_payload_uop_decoded_imm                           (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_imm[31:0]                    ), //o
    .io_commit_0_entry_payload_uop_decoded_immUsage                      (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_immUsage[2:0]                ), //o
    .io_commit_0_entry_payload_uop_decoded_aluCtrl_valid                 (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid                ), //o
    .io_commit_0_entry_payload_uop_decoded_aluCtrl_isSub                 (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_isSub                ), //o
    .io_commit_0_entry_payload_uop_decoded_aluCtrl_isAdd                 (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_isAdd                ), //o
    .io_commit_0_entry_payload_uop_decoded_aluCtrl_isSigned              (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_isSigned             ), //o
    .io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp[1:0]         ), //o
    .io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid              ), //o
    .io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRight             (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRight            ), //o
    .io_commit_0_entry_payload_uop_decoded_shiftCtrl_isArithmetic        (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_isArithmetic       ), //o
    .io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRotate            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRotate           ), //o
    .io_commit_0_entry_payload_uop_decoded_shiftCtrl_isDoubleWord        (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_shiftCtrl_isDoubleWord       ), //o
    .io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid              (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid             ), //o
    .io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isDiv              (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isDiv             ), //o
    .io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isSigned           (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isSigned          ), //o
    .io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isWordOp           (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isWordOp          ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_size                  (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_size[1:0]            ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad          (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad         ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_isStore               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isStore              ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_isLoadLinked          (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isLoadLinked         ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_isStoreCond           (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isStoreCond          ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_atomicOp              (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_atomicOp[4:0]        ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_isFence               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isFence              ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_fenceMode             (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_fenceMode[7:0]       ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_isCacheOp             (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isCacheOp            ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_cacheOpType           (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_cacheOpType[4:0]     ), //o
    .io_commit_0_entry_payload_uop_decoded_memCtrl_isPrefetch            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_memCtrl_isPrefetch           ), //o
    .io_commit_0_entry_payload_uop_decoded_branchCtrl_condition          (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition[4:0]    ), //o
    .io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump             (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump            ), //o
    .io_commit_0_entry_payload_uop_decoded_branchCtrl_isLink             (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_isLink            ), //o
    .io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx        (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx[4:0]  ), //o
    .io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype      (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype[1:0]), //o
    .io_commit_0_entry_payload_uop_decoded_branchCtrl_isIndirect         (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_isIndirect        ), //o
    .io_commit_0_entry_payload_uop_decoded_branchCtrl_laCfIdx            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchCtrl_laCfIdx[2:0]      ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[3:0]          ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1[1:0]      ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2[1:0]      ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest[1:0]      ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_roundingMode          (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_roundingMode[2:0]    ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_isIntegerDest         (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_isIntegerDest        ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_isSignedCvt           (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_isSignedCvt          ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_fmaNegSrc1            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fmaNegSrc1           ), //o
    .io_commit_0_entry_payload_uop_decoded_fpuCtrl_fcmpCond              (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fcmpCond[4:0]        ), //o
    .io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr[13:0]        ), //o
    .io_commit_0_entry_payload_uop_decoded_csrCtrl_isWrite               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_isWrite              ), //o
    .io_commit_0_entry_payload_uop_decoded_csrCtrl_isRead                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_isRead               ), //o
    .io_commit_0_entry_payload_uop_decoded_csrCtrl_isExchange            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_isExchange           ), //o
    .io_commit_0_entry_payload_uop_decoded_csrCtrl_useUimmAsSrc          (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_csrCtrl_useUimmAsSrc         ), //o
    .io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode[19:0]        ), //o
    .io_commit_0_entry_payload_uop_decoded_sysCtrl_isExceptionReturn     (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_sysCtrl_isExceptionReturn    ), //o
    .io_commit_0_entry_payload_uop_decoded_sysCtrl_isTlbOp               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_sysCtrl_isTlbOp              ), //o
    .io_commit_0_entry_payload_uop_decoded_sysCtrl_tlbOpType             (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_sysCtrl_tlbOpType[3:0]       ), //o
    .io_commit_0_entry_payload_uop_decoded_decodeExceptionCode           (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode[1:0]     ), //o
    .io_commit_0_entry_payload_uop_decoded_hasDecodeException            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_hasDecodeException           ), //o
    .io_commit_0_entry_payload_uop_decoded_isMicrocode                   (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isMicrocode                  ), //o
    .io_commit_0_entry_payload_uop_decoded_microcodeEntry                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_microcodeEntry[7:0]          ), //o
    .io_commit_0_entry_payload_uop_decoded_isSerializing                 (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isSerializing                ), //o
    .io_commit_0_entry_payload_uop_decoded_isBranchOrJump                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isBranchOrJump               ), //o
    .io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken      (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken     ), //o
    .io_commit_0_entry_payload_uop_decoded_branchPrediction_target       (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchPrediction_target[31:0]), //o
    .io_commit_0_entry_payload_uop_decoded_branchPrediction_wasPredicted (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_branchPrediction_wasPredicted), //o
    .io_commit_0_entry_payload_uop_rename_physSrc1_idx                   (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physSrc1_idx[5:0]             ), //o
    .io_commit_0_entry_payload_uop_rename_physSrc1IsFpr                  (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physSrc1IsFpr                 ), //o
    .io_commit_0_entry_payload_uop_rename_physSrc2_idx                   (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physSrc2_idx[5:0]             ), //o
    .io_commit_0_entry_payload_uop_rename_physSrc2IsFpr                  (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physSrc2IsFpr                 ), //o
    .io_commit_0_entry_payload_uop_rename_physDest_idx                   (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physDest_idx[5:0]             ), //o
    .io_commit_0_entry_payload_uop_rename_physDestIsFpr                  (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_physDestIsFpr                 ), //o
    .io_commit_0_entry_payload_uop_rename_oldPhysDest_idx                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_oldPhysDest_idx[5:0]          ), //o
    .io_commit_0_entry_payload_uop_rename_oldPhysDestIsFpr               (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_oldPhysDestIsFpr              ), //o
    .io_commit_0_entry_payload_uop_rename_allocatesPhysDest              (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_allocatesPhysDest             ), //o
    .io_commit_0_entry_payload_uop_rename_writesToPhysReg                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_writesToPhysReg               ), //o
    .io_commit_0_entry_payload_uop_robPtr                                (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_robPtr[3:0]                          ), //o
    .io_commit_0_entry_payload_uop_uniqueId                              (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_uniqueId[15:0]                       ), //o
    .io_commit_0_entry_payload_uop_dispatched                            (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_dispatched                           ), //o
    .io_commit_0_entry_payload_uop_executed                              (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_executed                             ), //o
    .io_commit_0_entry_payload_uop_hasException                          (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_hasException                         ), //o
    .io_commit_0_entry_payload_uop_exceptionCode                         (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_exceptionCode[7:0]                   ), //o
    .io_commit_0_entry_payload_pc                                        (ROBPlugin_robComponent_io_commit_0_entry_payload_pc[31:0]                                 ), //o
    .io_commit_0_entry_status_busy                                       (ROBPlugin_robComponent_io_commit_0_entry_status_busy                                      ), //o
    .io_commit_0_entry_status_done                                       (ROBPlugin_robComponent_io_commit_0_entry_status_done                                      ), //o
    .io_commit_0_entry_status_isMispredictedBranch                       (ROBPlugin_robComponent_io_commit_0_entry_status_isMispredictedBranch                      ), //o
    .io_commit_0_entry_status_isTaken                                    (ROBPlugin_robComponent_io_commit_0_entry_status_isTaken                                   ), //o
    .io_commit_0_entry_status_result                                     (ROBPlugin_robComponent_io_commit_0_entry_status_result[31:0]                              ), //o
    .io_commit_0_entry_status_hasException                               (ROBPlugin_robComponent_io_commit_0_entry_status_hasException                              ), //o
    .io_commit_0_entry_status_exceptionCode                              (ROBPlugin_robComponent_io_commit_0_entry_status_exceptionCode[7:0]                        ), //o
    .io_commit_0_entry_status_genBit                                     (ROBPlugin_robComponent_io_commit_0_entry_status_genBit                                    ), //o
    .io_commitAck_0                                                      (CommitPlugin_logic_s0_commitAckMasks_0                                                    ), //i
    .io_flush_valid                                                      (ROBPlugin_aggregatedFlushSignal_valid                                                     ), //i
    .io_flush_payload_reason                                             (ROBPlugin_aggregatedFlushSignal_payload_reason[1:0]                                       ), //i
    .io_flush_payload_targetRobPtr                                       (ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr[3:0]                                 ), //i
    .io_flushed                                                          (ROBPlugin_robComponent_io_flushed                                                         ), //o
    .io_empty                                                            (ROBPlugin_robComponent_io_empty                                                           ), //o
    .io_headPtrOut                                                       (ROBPlugin_robComponent_io_headPtrOut[3:0]                                                 ), //o
    .io_tailPtrOut                                                       (ROBPlugin_robComponent_io_tailPtrOut[3:0]                                                 ), //o
    .io_countOut                                                         (ROBPlugin_robComponent_io_countOut[3:0]                                                   ), //o
    .clk                                                                 (clk                                                                                       ), //i
    .reset                                                               (reset                                                                                     )  //i
  );
  RenameMapTable RenameMapTablePlugin_early_setup_rat (
    .io_readPorts_0_archReg                  (RenamePlugin_setup_renameUnit_io_ratReadPorts_0_archReg[4:0]                     ), //i
    .io_readPorts_0_physReg                  (RenameMapTablePlugin_early_setup_rat_io_readPorts_0_physReg[5:0]                 ), //o
    .io_readPorts_1_archReg                  (RenamePlugin_setup_renameUnit_io_ratReadPorts_1_archReg[4:0]                     ), //i
    .io_readPorts_1_physReg                  (RenameMapTablePlugin_early_setup_rat_io_readPorts_1_physReg[5:0]                 ), //o
    .io_readPorts_2_archReg                  (RenamePlugin_setup_renameUnit_io_ratReadPorts_2_archReg[4:0]                     ), //i
    .io_readPorts_2_physReg                  (RenameMapTablePlugin_early_setup_rat_io_readPorts_2_physReg[5:0]                 ), //o
    .io_writePorts_0_wen                     (RenameMapTablePlugin_early_setup_rat_io_writePorts_0_wen                         ), //i
    .io_writePorts_0_archReg                 (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archDest_idx[4:0]      ), //i
    .io_writePorts_0_physReg                 (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physDest_idx[5:0]       ), //i
    .io_currentState_mapping_0               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_0[5:0]              ), //o
    .io_currentState_mapping_1               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_1[5:0]              ), //o
    .io_currentState_mapping_2               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_2[5:0]              ), //o
    .io_currentState_mapping_3               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_3[5:0]              ), //o
    .io_currentState_mapping_4               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_4[5:0]              ), //o
    .io_currentState_mapping_5               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_5[5:0]              ), //o
    .io_currentState_mapping_6               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_6[5:0]              ), //o
    .io_currentState_mapping_7               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_7[5:0]              ), //o
    .io_currentState_mapping_8               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_8[5:0]              ), //o
    .io_currentState_mapping_9               (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_9[5:0]              ), //o
    .io_currentState_mapping_10              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_10[5:0]             ), //o
    .io_currentState_mapping_11              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_11[5:0]             ), //o
    .io_currentState_mapping_12              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_12[5:0]             ), //o
    .io_currentState_mapping_13              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_13[5:0]             ), //o
    .io_currentState_mapping_14              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_14[5:0]             ), //o
    .io_currentState_mapping_15              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_15[5:0]             ), //o
    .io_currentState_mapping_16              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_16[5:0]             ), //o
    .io_currentState_mapping_17              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_17[5:0]             ), //o
    .io_currentState_mapping_18              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_18[5:0]             ), //o
    .io_currentState_mapping_19              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_19[5:0]             ), //o
    .io_currentState_mapping_20              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_20[5:0]             ), //o
    .io_currentState_mapping_21              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_21[5:0]             ), //o
    .io_currentState_mapping_22              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_22[5:0]             ), //o
    .io_currentState_mapping_23              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_23[5:0]             ), //o
    .io_currentState_mapping_24              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_24[5:0]             ), //o
    .io_currentState_mapping_25              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_25[5:0]             ), //o
    .io_currentState_mapping_26              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_26[5:0]             ), //o
    .io_currentState_mapping_27              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_27[5:0]             ), //o
    .io_currentState_mapping_28              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_28[5:0]             ), //o
    .io_currentState_mapping_29              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_29[5:0]             ), //o
    .io_currentState_mapping_30              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_30[5:0]             ), //o
    .io_currentState_mapping_31              (RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_31[5:0]             ), //o
    .io_checkpointRestore_valid              (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_valid                  ), //i
    .io_checkpointRestore_ready              (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_ready                  ), //o
    .io_checkpointRestore_payload_mapping_0  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_0[5:0] ), //i
    .io_checkpointRestore_payload_mapping_1  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_1[5:0] ), //i
    .io_checkpointRestore_payload_mapping_2  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_2[5:0] ), //i
    .io_checkpointRestore_payload_mapping_3  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_3[5:0] ), //i
    .io_checkpointRestore_payload_mapping_4  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_4[5:0] ), //i
    .io_checkpointRestore_payload_mapping_5  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_5[5:0] ), //i
    .io_checkpointRestore_payload_mapping_6  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_6[5:0] ), //i
    .io_checkpointRestore_payload_mapping_7  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_7[5:0] ), //i
    .io_checkpointRestore_payload_mapping_8  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_8[5:0] ), //i
    .io_checkpointRestore_payload_mapping_9  (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_9[5:0] ), //i
    .io_checkpointRestore_payload_mapping_10 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_10[5:0]), //i
    .io_checkpointRestore_payload_mapping_11 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_11[5:0]), //i
    .io_checkpointRestore_payload_mapping_12 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_12[5:0]), //i
    .io_checkpointRestore_payload_mapping_13 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_13[5:0]), //i
    .io_checkpointRestore_payload_mapping_14 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_14[5:0]), //i
    .io_checkpointRestore_payload_mapping_15 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_15[5:0]), //i
    .io_checkpointRestore_payload_mapping_16 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_16[5:0]), //i
    .io_checkpointRestore_payload_mapping_17 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_17[5:0]), //i
    .io_checkpointRestore_payload_mapping_18 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_18[5:0]), //i
    .io_checkpointRestore_payload_mapping_19 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_19[5:0]), //i
    .io_checkpointRestore_payload_mapping_20 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_20[5:0]), //i
    .io_checkpointRestore_payload_mapping_21 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_21[5:0]), //i
    .io_checkpointRestore_payload_mapping_22 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_22[5:0]), //i
    .io_checkpointRestore_payload_mapping_23 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_23[5:0]), //i
    .io_checkpointRestore_payload_mapping_24 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_24[5:0]), //i
    .io_checkpointRestore_payload_mapping_25 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_25[5:0]), //i
    .io_checkpointRestore_payload_mapping_26 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_26[5:0]), //i
    .io_checkpointRestore_payload_mapping_27 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_27[5:0]), //i
    .io_checkpointRestore_payload_mapping_28 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_28[5:0]), //i
    .io_checkpointRestore_payload_mapping_29 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_29[5:0]), //i
    .io_checkpointRestore_payload_mapping_30 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_30[5:0]), //i
    .io_checkpointRestore_payload_mapping_31 (RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_31[5:0]), //i
    .io_checkpointSave_valid                 (                                                                                 ), //i
    .io_checkpointSave_ready                 (RenameMapTablePlugin_early_setup_rat_io_checkpointSave_ready                     ), //o
    .io_checkpointSave_payload_mapping_0     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_1     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_2     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_3     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_4     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_5     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_6     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_7     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_8     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_9     (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_10    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_11    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_12    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_13    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_14    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_15    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_16    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_17    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_18    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_19    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_20    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_21    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_22    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_23    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_24    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_25    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_26    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_27    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_28    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_29    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_30    (                                                                                 ), //i
    .io_checkpointSave_payload_mapping_31    (                                                                                 ), //i
    .clk                                     (clk                                                                              ), //i
    .reset                                   (reset                                                                            )  //i
  );
  SimpleFreeList SimpleFreeListPlugin_early_setup_freeList (
    .io_allocate_0_enable  (SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_enable                  ), //i
    .io_allocate_0_physReg (SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_physReg[5:0]            ), //o
    .io_allocate_0_success (SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_success                 ), //o
    .io_free_0_enable      (when_CommitPlugin_l265                                                          ), //i
    .io_free_0_physReg     (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_oldPhysDest_idx[5:0]), //i
    .io_recover            (SimpleFreeListPlugin_early_setup_freeList_io_recover                            ), //i
    .io_numFreeRegs        (SimpleFreeListPlugin_early_setup_freeList_io_numFreeRegs[5:0]                   ), //o
    .clk                   (clk                                                                             ), //i
    .reset                 (reset                                                                           )  //i
  );
  OneShot oneShot_14 (
    .io_triggerIn (oneShot_14_io_triggerIn), //i
    .io_pulseOut  (oneShot_14_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  OneShot oneShot_15 (
    .io_triggerIn (oneShot_15_io_triggerIn), //i
    .io_pulseOut  (oneShot_15_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  OneShot oneShot_16 (
    .io_triggerIn (oneShot_16_io_triggerIn), //i
    .io_pulseOut  (oneShot_16_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  OneShot oneShot_17 (
    .io_triggerIn (oneShot_17_io_triggerIn), //i
    .io_pulseOut  (oneShot_17_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  RenameUnit RenamePlugin_setup_renameUnit (
    .io_decodedUopsIn_0_pc                                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_pc[31:0]                               ), //i
    .io_decodedUopsIn_0_isValid                                (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isValid                                ), //i
    .io_decodedUopsIn_0_uopCode                                (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode[4:0]                           ), //i
    .io_decodedUopsIn_0_exeUnit                                (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit[3:0]                           ), //i
    .io_decodedUopsIn_0_isa                                    (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa[1:0]                               ), //i
    .io_decodedUopsIn_0_archDest_idx                           (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx[4:0]                      ), //i
    .io_decodedUopsIn_0_archDest_rtype                         (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype[1:0]                    ), //i
    .io_decodedUopsIn_0_writeArchDestEn                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn                        ), //i
    .io_decodedUopsIn_0_archSrc1_idx                           (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx[4:0]                      ), //i
    .io_decodedUopsIn_0_archSrc1_rtype                         (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype[1:0]                    ), //i
    .io_decodedUopsIn_0_useArchSrc1                            (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1                            ), //i
    .io_decodedUopsIn_0_archSrc2_idx                           (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx[4:0]                      ), //i
    .io_decodedUopsIn_0_archSrc2_rtype                         (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype[1:0]                    ), //i
    .io_decodedUopsIn_0_useArchSrc2                            (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2                            ), //i
    .io_decodedUopsIn_0_usePcForAddr                           (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr                           ), //i
    .io_decodedUopsIn_0_imm                                    (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_imm[31:0]                              ), //i
    .io_decodedUopsIn_0_immUsage                               (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage[2:0]                          ), //i
    .io_decodedUopsIn_0_aluCtrl_valid                          (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid                          ), //i
    .io_decodedUopsIn_0_aluCtrl_isSub                          (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub                          ), //i
    .io_decodedUopsIn_0_aluCtrl_isAdd                          (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd                          ), //i
    .io_decodedUopsIn_0_aluCtrl_isSigned                       (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned                       ), //i
    .io_decodedUopsIn_0_aluCtrl_logicOp                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp[1:0]                   ), //i
    .io_decodedUopsIn_0_shiftCtrl_valid                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid                        ), //i
    .io_decodedUopsIn_0_shiftCtrl_isRight                      (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight                      ), //i
    .io_decodedUopsIn_0_shiftCtrl_isArithmetic                 (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic                 ), //i
    .io_decodedUopsIn_0_shiftCtrl_isRotate                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate                     ), //i
    .io_decodedUopsIn_0_shiftCtrl_isDoubleWord                 (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord                 ), //i
    .io_decodedUopsIn_0_mulDivCtrl_valid                       (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid                       ), //i
    .io_decodedUopsIn_0_mulDivCtrl_isDiv                       (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv                       ), //i
    .io_decodedUopsIn_0_mulDivCtrl_isSigned                    (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned                    ), //i
    .io_decodedUopsIn_0_mulDivCtrl_isWordOp                    (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp                    ), //i
    .io_decodedUopsIn_0_memCtrl_size                           (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size[1:0]                      ), //i
    .io_decodedUopsIn_0_memCtrl_isSignedLoad                   (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad                   ), //i
    .io_decodedUopsIn_0_memCtrl_isStore                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore                        ), //i
    .io_decodedUopsIn_0_memCtrl_isLoadLinked                   (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked                   ), //i
    .io_decodedUopsIn_0_memCtrl_isStoreCond                    (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond                    ), //i
    .io_decodedUopsIn_0_memCtrl_atomicOp                       (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp[4:0]                  ), //i
    .io_decodedUopsIn_0_memCtrl_isFence                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence                        ), //i
    .io_decodedUopsIn_0_memCtrl_fenceMode                      (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode[7:0]                 ), //i
    .io_decodedUopsIn_0_memCtrl_isCacheOp                      (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp                      ), //i
    .io_decodedUopsIn_0_memCtrl_cacheOpType                    (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType[4:0]               ), //i
    .io_decodedUopsIn_0_memCtrl_isPrefetch                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch                     ), //i
    .io_decodedUopsIn_0_branchCtrl_condition                   (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition[4:0]              ), //i
    .io_decodedUopsIn_0_branchCtrl_isJump                      (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump                      ), //i
    .io_decodedUopsIn_0_branchCtrl_isLink                      (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink                      ), //i
    .io_decodedUopsIn_0_branchCtrl_linkReg_idx                 (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx[4:0]            ), //i
    .io_decodedUopsIn_0_branchCtrl_linkReg_rtype               (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype[1:0]          ), //i
    .io_decodedUopsIn_0_branchCtrl_isIndirect                  (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect                  ), //i
    .io_decodedUopsIn_0_branchCtrl_laCfIdx                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx[2:0]                ), //i
    .io_decodedUopsIn_0_fpuCtrl_opType                         (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType[3:0]                    ), //i
    .io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1[1:0]                ), //i
    .io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2[1:0]                ), //i
    .io_decodedUopsIn_0_fpuCtrl_fpSizeDest                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest[1:0]                ), //i
    .io_decodedUopsIn_0_fpuCtrl_roundingMode                   (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode[2:0]              ), //i
    .io_decodedUopsIn_0_fpuCtrl_isIntegerDest                  (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest                  ), //i
    .io_decodedUopsIn_0_fpuCtrl_isSignedCvt                    (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt                    ), //i
    .io_decodedUopsIn_0_fpuCtrl_fmaNegSrc1                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1                     ), //i
    .io_decodedUopsIn_0_fpuCtrl_fcmpCond                       (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond[4:0]                  ), //i
    .io_decodedUopsIn_0_csrCtrl_csrAddr                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr[13:0]                  ), //i
    .io_decodedUopsIn_0_csrCtrl_isWrite                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite                        ), //i
    .io_decodedUopsIn_0_csrCtrl_isRead                         (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead                         ), //i
    .io_decodedUopsIn_0_csrCtrl_isExchange                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange                     ), //i
    .io_decodedUopsIn_0_csrCtrl_useUimmAsSrc                   (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc                   ), //i
    .io_decodedUopsIn_0_sysCtrl_sysCode                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode[19:0]                  ), //i
    .io_decodedUopsIn_0_sysCtrl_isExceptionReturn              (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn              ), //i
    .io_decodedUopsIn_0_sysCtrl_isTlbOp                        (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp                        ), //i
    .io_decodedUopsIn_0_sysCtrl_tlbOpType                      (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType[3:0]                 ), //i
    .io_decodedUopsIn_0_decodeExceptionCode                    (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode[1:0]               ), //i
    .io_decodedUopsIn_0_hasDecodeException                     (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException                     ), //i
    .io_decodedUopsIn_0_isMicrocode                            (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode                            ), //i
    .io_decodedUopsIn_0_microcodeEntry                         (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry[7:0]                    ), //i
    .io_decodedUopsIn_0_isSerializing                          (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isSerializing                          ), //i
    .io_decodedUopsIn_0_isBranchOrJump                         (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump                         ), //i
    .io_decodedUopsIn_0_branchPrediction_isTaken               (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken               ), //i
    .io_decodedUopsIn_0_branchPrediction_target                (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target[31:0]          ), //i
    .io_decodedUopsIn_0_branchPrediction_wasPredicted          (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted          ), //i
    .io_physRegsIn_0                                           (SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_physReg[5:0]                   ), //i
    .io_renamedUopsOut_0_decoded_pc                            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_pc[31:0]                     ), //o
    .io_renamedUopsOut_0_decoded_isValid                       (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isValid                      ), //o
    .io_renamedUopsOut_0_decoded_uopCode                       (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_uopCode[4:0]                 ), //o
    .io_renamedUopsOut_0_decoded_exeUnit                       (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_exeUnit[3:0]                 ), //o
    .io_renamedUopsOut_0_decoded_isa                           (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isa[1:0]                     ), //o
    .io_renamedUopsOut_0_decoded_archDest_idx                  (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archDest_idx[4:0]            ), //o
    .io_renamedUopsOut_0_decoded_archDest_rtype                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archDest_rtype[1:0]          ), //o
    .io_renamedUopsOut_0_decoded_writeArchDestEn               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_writeArchDestEn              ), //o
    .io_renamedUopsOut_0_decoded_archSrc1_idx                  (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc1_idx[4:0]            ), //o
    .io_renamedUopsOut_0_decoded_archSrc1_rtype                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc1_rtype[1:0]          ), //o
    .io_renamedUopsOut_0_decoded_useArchSrc1                   (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_useArchSrc1                  ), //o
    .io_renamedUopsOut_0_decoded_archSrc2_idx                  (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc2_idx[4:0]            ), //o
    .io_renamedUopsOut_0_decoded_archSrc2_rtype                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc2_rtype[1:0]          ), //o
    .io_renamedUopsOut_0_decoded_useArchSrc2                   (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_useArchSrc2                  ), //o
    .io_renamedUopsOut_0_decoded_usePcForAddr                  (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_usePcForAddr                 ), //o
    .io_renamedUopsOut_0_decoded_imm                           (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_imm[31:0]                    ), //o
    .io_renamedUopsOut_0_decoded_immUsage                      (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_immUsage[2:0]                ), //o
    .io_renamedUopsOut_0_decoded_aluCtrl_valid                 (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_valid                ), //o
    .io_renamedUopsOut_0_decoded_aluCtrl_isSub                 (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isSub                ), //o
    .io_renamedUopsOut_0_decoded_aluCtrl_isAdd                 (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isAdd                ), //o
    .io_renamedUopsOut_0_decoded_aluCtrl_isSigned              (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isSigned             ), //o
    .io_renamedUopsOut_0_decoded_aluCtrl_logicOp               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_logicOp[1:0]         ), //o
    .io_renamedUopsOut_0_decoded_shiftCtrl_valid               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_valid              ), //o
    .io_renamedUopsOut_0_decoded_shiftCtrl_isRight             (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isRight            ), //o
    .io_renamedUopsOut_0_decoded_shiftCtrl_isArithmetic        (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isArithmetic       ), //o
    .io_renamedUopsOut_0_decoded_shiftCtrl_isRotate            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isRotate           ), //o
    .io_renamedUopsOut_0_decoded_shiftCtrl_isDoubleWord        (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isDoubleWord       ), //o
    .io_renamedUopsOut_0_decoded_mulDivCtrl_valid              (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_valid             ), //o
    .io_renamedUopsOut_0_decoded_mulDivCtrl_isDiv              (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isDiv             ), //o
    .io_renamedUopsOut_0_decoded_mulDivCtrl_isSigned           (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isSigned          ), //o
    .io_renamedUopsOut_0_decoded_mulDivCtrl_isWordOp           (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isWordOp          ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_size                  (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_size[1:0]            ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_isSignedLoad          (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isSignedLoad         ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_isStore               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isStore              ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_isLoadLinked          (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isLoadLinked         ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_isStoreCond           (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isStoreCond          ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_atomicOp              (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_atomicOp[4:0]        ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_isFence               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isFence              ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_fenceMode             (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_fenceMode[7:0]       ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_isCacheOp             (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isCacheOp            ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_cacheOpType           (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_cacheOpType[4:0]     ), //o
    .io_renamedUopsOut_0_decoded_memCtrl_isPrefetch            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isPrefetch           ), //o
    .io_renamedUopsOut_0_decoded_branchCtrl_condition          (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_condition[4:0]    ), //o
    .io_renamedUopsOut_0_decoded_branchCtrl_isJump             (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isJump            ), //o
    .io_renamedUopsOut_0_decoded_branchCtrl_isLink             (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isLink            ), //o
    .io_renamedUopsOut_0_decoded_branchCtrl_linkReg_idx        (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_linkReg_idx[4:0]  ), //o
    .io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype      (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype[1:0]), //o
    .io_renamedUopsOut_0_decoded_branchCtrl_isIndirect         (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isIndirect        ), //o
    .io_renamedUopsOut_0_decoded_branchCtrl_laCfIdx            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_laCfIdx[2:0]      ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_opType                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_opType[3:0]          ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1[1:0]      ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2[1:0]      ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest[1:0]      ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_roundingMode          (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_roundingMode[2:0]    ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_isIntegerDest         (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_isIntegerDest        ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_isSignedCvt           (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_isSignedCvt          ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_fmaNegSrc1            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fmaNegSrc1           ), //o
    .io_renamedUopsOut_0_decoded_fpuCtrl_fcmpCond              (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fcmpCond[4:0]        ), //o
    .io_renamedUopsOut_0_decoded_csrCtrl_csrAddr               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_csrAddr[13:0]        ), //o
    .io_renamedUopsOut_0_decoded_csrCtrl_isWrite               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isWrite              ), //o
    .io_renamedUopsOut_0_decoded_csrCtrl_isRead                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isRead               ), //o
    .io_renamedUopsOut_0_decoded_csrCtrl_isExchange            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isExchange           ), //o
    .io_renamedUopsOut_0_decoded_csrCtrl_useUimmAsSrc          (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_useUimmAsSrc         ), //o
    .io_renamedUopsOut_0_decoded_sysCtrl_sysCode               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_sysCode[19:0]        ), //o
    .io_renamedUopsOut_0_decoded_sysCtrl_isExceptionReturn     (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_isExceptionReturn    ), //o
    .io_renamedUopsOut_0_decoded_sysCtrl_isTlbOp               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_isTlbOp              ), //o
    .io_renamedUopsOut_0_decoded_sysCtrl_tlbOpType             (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_tlbOpType[3:0]       ), //o
    .io_renamedUopsOut_0_decoded_decodeExceptionCode           (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_decodeExceptionCode[1:0]     ), //o
    .io_renamedUopsOut_0_decoded_hasDecodeException            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_hasDecodeException           ), //o
    .io_renamedUopsOut_0_decoded_isMicrocode                   (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isMicrocode                  ), //o
    .io_renamedUopsOut_0_decoded_microcodeEntry                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_microcodeEntry[7:0]          ), //o
    .io_renamedUopsOut_0_decoded_isSerializing                 (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isSerializing                ), //o
    .io_renamedUopsOut_0_decoded_isBranchOrJump                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isBranchOrJump               ), //o
    .io_renamedUopsOut_0_decoded_branchPrediction_isTaken      (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_isTaken     ), //o
    .io_renamedUopsOut_0_decoded_branchPrediction_target       (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_target[31:0]), //o
    .io_renamedUopsOut_0_decoded_branchPrediction_wasPredicted (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_wasPredicted), //o
    .io_renamedUopsOut_0_rename_physSrc1_idx                   (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc1_idx[5:0]             ), //o
    .io_renamedUopsOut_0_rename_physSrc1IsFpr                  (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc1IsFpr                 ), //o
    .io_renamedUopsOut_0_rename_physSrc2_idx                   (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc2_idx[5:0]             ), //o
    .io_renamedUopsOut_0_rename_physSrc2IsFpr                  (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc2IsFpr                 ), //o
    .io_renamedUopsOut_0_rename_physDest_idx                   (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physDest_idx[5:0]             ), //o
    .io_renamedUopsOut_0_rename_physDestIsFpr                  (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physDestIsFpr                 ), //o
    .io_renamedUopsOut_0_rename_oldPhysDest_idx                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_oldPhysDest_idx[5:0]          ), //o
    .io_renamedUopsOut_0_rename_oldPhysDestIsFpr               (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_oldPhysDestIsFpr              ), //o
    .io_renamedUopsOut_0_rename_allocatesPhysDest              (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_allocatesPhysDest             ), //o
    .io_renamedUopsOut_0_rename_writesToPhysReg                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_writesToPhysReg               ), //o
    .io_renamedUopsOut_0_robPtr                                (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_robPtr[3:0]                          ), //o
    .io_renamedUopsOut_0_uniqueId                              (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_uniqueId[15:0]                       ), //o
    .io_renamedUopsOut_0_dispatched                            (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_dispatched                           ), //o
    .io_renamedUopsOut_0_executed                              (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_executed                             ), //o
    .io_renamedUopsOut_0_hasException                          (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_hasException                         ), //o
    .io_renamedUopsOut_0_exceptionCode                         (RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_exceptionCode[7:0]                   ), //o
    .io_numPhysRegsRequired                                    (RenamePlugin_setup_renameUnit_io_numPhysRegsRequired                                   ), //o
    .io_ratReadPorts_0_archReg                                 (RenamePlugin_setup_renameUnit_io_ratReadPorts_0_archReg[4:0]                           ), //o
    .io_ratReadPorts_0_physReg                                 (RenameMapTablePlugin_early_setup_rat_io_readPorts_0_physReg[5:0]                       ), //i
    .io_ratReadPorts_1_archReg                                 (RenamePlugin_setup_renameUnit_io_ratReadPorts_1_archReg[4:0]                           ), //o
    .io_ratReadPorts_1_physReg                                 (RenameMapTablePlugin_early_setup_rat_io_readPorts_1_physReg[5:0]                       ), //i
    .io_ratReadPorts_2_archReg                                 (RenamePlugin_setup_renameUnit_io_ratReadPorts_2_archReg[4:0]                           ), //o
    .io_ratReadPorts_2_physReg                                 (RenameMapTablePlugin_early_setup_rat_io_readPorts_2_physReg[5:0]                       ), //i
    .io_ratWritePorts_0_wen                                    (RenamePlugin_setup_renameUnit_io_ratWritePorts_0_wen                                   ), //o
    .io_ratWritePorts_0_archReg                                (RenamePlugin_setup_renameUnit_io_ratWritePorts_0_archReg[4:0]                          ), //o
    .io_ratWritePorts_0_physReg                                (RenamePlugin_setup_renameUnit_io_ratWritePorts_0_physReg[5:0]                          ), //o
    .clk                                                       (clk                                                                                    ), //i
    .reset                                                     (reset                                                                                  )  //i
  );
  EightSegmentDisplayController DebugDisplayPlugin_hw_dpyController (
    .io_value    (_zz_when_Debug_l71[7:0]                             ), //i
    .io_dp0      (DebugDisplayPlugin_hw_dpyController_io_dp0          ), //i
    .io_dp1      (DebugDisplayPlugin_logic_displayArea_dpToggle       ), //i
    .io_dpy0_out (DebugDisplayPlugin_hw_dpyController_io_dpy0_out[7:0]), //o
    .io_dpy1_out (DebugDisplayPlugin_hw_dpyController_io_dpy1_out[7:0])  //o
  );
  StreamArbiter_6 streamArbiter_8 (
    .io_inputs_0_valid                 (AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_valid                     ), //i
    .io_inputs_0_ready                 (streamArbiter_8_io_inputs_0_ready                                           ), //o
    .io_inputs_0_payload_physRegIdx    (AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_physRegIdx[5:0]   ), //i
    .io_inputs_0_payload_physRegData   (AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_physRegData[31:0] ), //i
    .io_inputs_0_payload_robPtr        (AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_robPtr[3:0]       ), //i
    .io_inputs_0_payload_isFPR         (AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_isFPR             ), //i
    .io_inputs_0_payload_hasException  (AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_hasException      ), //i
    .io_inputs_0_payload_exceptionCode (AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_exceptionCode[7:0]), //i
    .io_inputs_1_valid                 (MulEU_MulEuPlugin_bypassOutputPort_toStream_valid                           ), //i
    .io_inputs_1_ready                 (streamArbiter_8_io_inputs_1_ready                                           ), //o
    .io_inputs_1_payload_physRegIdx    (MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_physRegIdx[5:0]         ), //i
    .io_inputs_1_payload_physRegData   (MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_physRegData[31:0]       ), //i
    .io_inputs_1_payload_robPtr        (MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_robPtr[3:0]             ), //i
    .io_inputs_1_payload_isFPR         (MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_isFPR                   ), //i
    .io_inputs_1_payload_hasException  (MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_hasException            ), //i
    .io_inputs_1_payload_exceptionCode (MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_exceptionCode[7:0]      ), //i
    .io_inputs_2_valid                 (BranchEU_BranchEuPlugin_bypassOutputPort_toStream_valid                     ), //i
    .io_inputs_2_ready                 (streamArbiter_8_io_inputs_2_ready                                           ), //o
    .io_inputs_2_payload_physRegIdx    (BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_physRegIdx[5:0]   ), //i
    .io_inputs_2_payload_physRegData   (BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_physRegData[31:0] ), //i
    .io_inputs_2_payload_robPtr        (BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_robPtr[3:0]       ), //i
    .io_inputs_2_payload_isFPR         (BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_isFPR             ), //i
    .io_inputs_2_payload_hasException  (BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_hasException      ), //i
    .io_inputs_2_payload_exceptionCode (BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_exceptionCode[7:0]), //i
    .io_output_valid                   (streamArbiter_8_io_output_valid                                             ), //o
    .io_output_ready                   (io_output_combStage_ready                                                   ), //i
    .io_output_payload_physRegIdx      (streamArbiter_8_io_output_payload_physRegIdx[5:0]                           ), //o
    .io_output_payload_physRegData     (streamArbiter_8_io_output_payload_physRegData[31:0]                         ), //o
    .io_output_payload_robPtr          (streamArbiter_8_io_output_payload_robPtr[3:0]                               ), //o
    .io_output_payload_isFPR           (streamArbiter_8_io_output_payload_isFPR                                     ), //o
    .io_output_payload_hasException    (streamArbiter_8_io_output_payload_hasException                              ), //o
    .io_output_payload_exceptionCode   (streamArbiter_8_io_output_payload_exceptionCode[7:0]                        ), //o
    .io_chosen                         (streamArbiter_8_io_chosen[1:0]                                              ), //o
    .io_chosenOH                       (streamArbiter_8_io_chosenOH[2:0]                                            ), //o
    .clk                               (clk                                                                         ), //i
    .reset                             (reset                                                                       )  //i
  );
  OneShot oneShot_18 (
    .io_triggerIn (oneShot_18_io_triggerIn), //i
    .io_pulseOut  (oneShot_18_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  OneShot oneShot_19 (
    .io_triggerIn (CommitPlugin_commitOOBReg), //i
    .io_pulseOut  (oneShot_19_io_pulseOut   ), //o
    .clk          (clk                      ), //i
    .reset        (reset                    )  //i
  );
  LA32RSimpleDecoder lA32RSimpleDecoder_1 (
    .io_instruction                              (s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_0[31:0]      ), //i
    .io_pcIn                                     (lA32RSimpleDecoder_1_io_pcIn[31:0]                              ), //i
    .io_decodedUop_pc                            (lA32RSimpleDecoder_1_io_decodedUop_pc[31:0]                     ), //o
    .io_decodedUop_isValid                       (lA32RSimpleDecoder_1_io_decodedUop_isValid                      ), //o
    .io_decodedUop_uopCode                       (lA32RSimpleDecoder_1_io_decodedUop_uopCode[4:0]                 ), //o
    .io_decodedUop_exeUnit                       (lA32RSimpleDecoder_1_io_decodedUop_exeUnit[3:0]                 ), //o
    .io_decodedUop_isa                           (lA32RSimpleDecoder_1_io_decodedUop_isa[1:0]                     ), //o
    .io_decodedUop_archDest_idx                  (lA32RSimpleDecoder_1_io_decodedUop_archDest_idx[4:0]            ), //o
    .io_decodedUop_archDest_rtype                (lA32RSimpleDecoder_1_io_decodedUop_archDest_rtype[1:0]          ), //o
    .io_decodedUop_writeArchDestEn               (lA32RSimpleDecoder_1_io_decodedUop_writeArchDestEn              ), //o
    .io_decodedUop_archSrc1_idx                  (lA32RSimpleDecoder_1_io_decodedUop_archSrc1_idx[4:0]            ), //o
    .io_decodedUop_archSrc1_rtype                (lA32RSimpleDecoder_1_io_decodedUop_archSrc1_rtype[1:0]          ), //o
    .io_decodedUop_useArchSrc1                   (lA32RSimpleDecoder_1_io_decodedUop_useArchSrc1                  ), //o
    .io_decodedUop_archSrc2_idx                  (lA32RSimpleDecoder_1_io_decodedUop_archSrc2_idx[4:0]            ), //o
    .io_decodedUop_archSrc2_rtype                (lA32RSimpleDecoder_1_io_decodedUop_archSrc2_rtype[1:0]          ), //o
    .io_decodedUop_useArchSrc2                   (lA32RSimpleDecoder_1_io_decodedUop_useArchSrc2                  ), //o
    .io_decodedUop_usePcForAddr                  (lA32RSimpleDecoder_1_io_decodedUop_usePcForAddr                 ), //o
    .io_decodedUop_imm                           (lA32RSimpleDecoder_1_io_decodedUop_imm[31:0]                    ), //o
    .io_decodedUop_immUsage                      (lA32RSimpleDecoder_1_io_decodedUop_immUsage[2:0]                ), //o
    .io_decodedUop_aluCtrl_valid                 (lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_valid                ), //o
    .io_decodedUop_aluCtrl_isSub                 (lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isSub                ), //o
    .io_decodedUop_aluCtrl_isAdd                 (lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isAdd                ), //o
    .io_decodedUop_aluCtrl_isSigned              (lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isSigned             ), //o
    .io_decodedUop_aluCtrl_logicOp               (lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_logicOp[1:0]         ), //o
    .io_decodedUop_shiftCtrl_valid               (lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_valid              ), //o
    .io_decodedUop_shiftCtrl_isRight             (lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isRight            ), //o
    .io_decodedUop_shiftCtrl_isArithmetic        (lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isArithmetic       ), //o
    .io_decodedUop_shiftCtrl_isRotate            (lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isRotate           ), //o
    .io_decodedUop_shiftCtrl_isDoubleWord        (lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isDoubleWord       ), //o
    .io_decodedUop_mulDivCtrl_valid              (lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_valid             ), //o
    .io_decodedUop_mulDivCtrl_isDiv              (lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isDiv             ), //o
    .io_decodedUop_mulDivCtrl_isSigned           (lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isSigned          ), //o
    .io_decodedUop_mulDivCtrl_isWordOp           (lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isWordOp          ), //o
    .io_decodedUop_memCtrl_size                  (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_size[1:0]            ), //o
    .io_decodedUop_memCtrl_isSignedLoad          (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isSignedLoad         ), //o
    .io_decodedUop_memCtrl_isStore               (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isStore              ), //o
    .io_decodedUop_memCtrl_isLoadLinked          (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isLoadLinked         ), //o
    .io_decodedUop_memCtrl_isStoreCond           (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isStoreCond          ), //o
    .io_decodedUop_memCtrl_atomicOp              (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_atomicOp[4:0]        ), //o
    .io_decodedUop_memCtrl_isFence               (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isFence              ), //o
    .io_decodedUop_memCtrl_fenceMode             (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_fenceMode[7:0]       ), //o
    .io_decodedUop_memCtrl_isCacheOp             (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isCacheOp            ), //o
    .io_decodedUop_memCtrl_cacheOpType           (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_cacheOpType[4:0]     ), //o
    .io_decodedUop_memCtrl_isPrefetch            (lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isPrefetch           ), //o
    .io_decodedUop_branchCtrl_condition          (lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_condition[4:0]    ), //o
    .io_decodedUop_branchCtrl_isJump             (lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isJump            ), //o
    .io_decodedUop_branchCtrl_isLink             (lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isLink            ), //o
    .io_decodedUop_branchCtrl_linkReg_idx        (lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_linkReg_idx[4:0]  ), //o
    .io_decodedUop_branchCtrl_linkReg_rtype      (lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_linkReg_rtype[1:0]), //o
    .io_decodedUop_branchCtrl_isIndirect         (lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isIndirect        ), //o
    .io_decodedUop_branchCtrl_laCfIdx            (lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_laCfIdx[2:0]      ), //o
    .io_decodedUop_fpuCtrl_opType                (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_opType[3:0]          ), //o
    .io_decodedUop_fpuCtrl_fpSizeSrc1            (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeSrc1[1:0]      ), //o
    .io_decodedUop_fpuCtrl_fpSizeSrc2            (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeSrc2[1:0]      ), //o
    .io_decodedUop_fpuCtrl_fpSizeDest            (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeDest[1:0]      ), //o
    .io_decodedUop_fpuCtrl_roundingMode          (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_roundingMode[2:0]    ), //o
    .io_decodedUop_fpuCtrl_isIntegerDest         (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_isIntegerDest        ), //o
    .io_decodedUop_fpuCtrl_isSignedCvt           (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_isSignedCvt          ), //o
    .io_decodedUop_fpuCtrl_fmaNegSrc1            (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fmaNegSrc1           ), //o
    .io_decodedUop_fpuCtrl_fcmpCond              (lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fcmpCond[4:0]        ), //o
    .io_decodedUop_csrCtrl_csrAddr               (lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_csrAddr[13:0]        ), //o
    .io_decodedUop_csrCtrl_isWrite               (lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isWrite              ), //o
    .io_decodedUop_csrCtrl_isRead                (lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isRead               ), //o
    .io_decodedUop_csrCtrl_isExchange            (lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isExchange           ), //o
    .io_decodedUop_csrCtrl_useUimmAsSrc          (lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_useUimmAsSrc         ), //o
    .io_decodedUop_sysCtrl_sysCode               (lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_sysCode[19:0]        ), //o
    .io_decodedUop_sysCtrl_isExceptionReturn     (lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_isExceptionReturn    ), //o
    .io_decodedUop_sysCtrl_isTlbOp               (lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_isTlbOp              ), //o
    .io_decodedUop_sysCtrl_tlbOpType             (lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_tlbOpType[3:0]       ), //o
    .io_decodedUop_decodeExceptionCode           (lA32RSimpleDecoder_1_io_decodedUop_decodeExceptionCode[1:0]     ), //o
    .io_decodedUop_hasDecodeException            (lA32RSimpleDecoder_1_io_decodedUop_hasDecodeException           ), //o
    .io_decodedUop_isMicrocode                   (lA32RSimpleDecoder_1_io_decodedUop_isMicrocode                  ), //o
    .io_decodedUop_microcodeEntry                (lA32RSimpleDecoder_1_io_decodedUop_microcodeEntry[7:0]          ), //o
    .io_decodedUop_isSerializing                 (lA32RSimpleDecoder_1_io_decodedUop_isSerializing                ), //o
    .io_decodedUop_isBranchOrJump                (lA32RSimpleDecoder_1_io_decodedUop_isBranchOrJump               ), //o
    .io_decodedUop_branchPrediction_isTaken      (lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_isTaken     ), //o
    .io_decodedUop_branchPrediction_target       (lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_target[31:0]), //o
    .io_decodedUop_branchPrediction_wasPredicted (lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_wasPredicted)  //o
  );
  IssueQueueComponent issueQueueComponent_4 (
    .io_allocateIn_valid                                             (DispatchPlugin_logic_iqRegs_0_1_valid                                            ), //i
    .io_allocateIn_ready                                             (issueQueueComponent_4_io_allocateIn_ready                                        ), //o
    .io_allocateIn_payload_uop_decoded_pc                            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_pc[31:0]                     ), //i
    .io_allocateIn_payload_uop_decoded_isValid                       (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isValid                      ), //i
    .io_allocateIn_payload_uop_decoded_uopCode                       (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode[4:0]                 ), //i
    .io_allocateIn_payload_uop_decoded_exeUnit                       (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit[3:0]                 ), //i
    .io_allocateIn_payload_uop_decoded_isa                           (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa[1:0]                     ), //i
    .io_allocateIn_payload_uop_decoded_archDest_idx                  (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archDest_rtype                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_writeArchDestEn               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_writeArchDestEn              ), //i
    .io_allocateIn_payload_uop_decoded_archSrc1_idx                  (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archSrc1_rtype                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_useArchSrc1                   (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_useArchSrc1                  ), //i
    .io_allocateIn_payload_uop_decoded_archSrc2_idx                  (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archSrc2_rtype                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_useArchSrc2                   (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_useArchSrc2                  ), //i
    .io_allocateIn_payload_uop_decoded_usePcForAddr                  (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_usePcForAddr                 ), //i
    .io_allocateIn_payload_uop_decoded_imm                           (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_imm[31:0]                    ), //i
    .io_allocateIn_payload_uop_decoded_immUsage                      (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage[2:0]                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_valid                 (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_valid                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isSub                 (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isSub                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isAdd                 (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isAdd                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isSigned              (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isSigned             ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_logicOp               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp[1:0]         ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_valid               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_valid              ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isRight             (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isRight            ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic        (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isArithmetic       ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isRotate           ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord        (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isDoubleWord       ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_valid              (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_valid             ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv              (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isDiv             ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned           (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isSigned          ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp           (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isWordOp          ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_size                  (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size[1:0]            ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad          (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isSignedLoad         ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isStore               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isStore              ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked          (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isLoadLinked         ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond           (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isStoreCond          ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_atomicOp              (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_atomicOp[4:0]        ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isFence               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isFence              ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_fenceMode             (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_fenceMode[7:0]       ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp             (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isCacheOp            ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType           (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_cacheOpType[4:0]     ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isPrefetch           ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_condition          (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition[4:0]    ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isJump             (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isJump            ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isLink             (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isLink            ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx        (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_idx[4:0]  ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype      (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype[1:0]), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect         (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isIndirect        ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_laCfIdx[2:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_opType                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_opType[3:0]          ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode          (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_roundingMode[2:0]    ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest         (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_isIntegerDest        ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt           (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_isSignedCvt          ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1           ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond              (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fcmpCond[4:0]        ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_csrAddr[13:0]        ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isWrite               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isWrite              ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isRead                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isRead               ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isExchange            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isExchange           ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc          (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_useUimmAsSrc         ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_sysCode               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_sysCode[19:0]        ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn     (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_isExceptionReturn    ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_isTlbOp              ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType             (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_tlbOpType[3:0]       ), //i
    .io_allocateIn_payload_uop_decoded_decodeExceptionCode           (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode[1:0]     ), //i
    .io_allocateIn_payload_uop_decoded_hasDecodeException            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_hasDecodeException           ), //i
    .io_allocateIn_payload_uop_decoded_isMicrocode                   (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isMicrocode                  ), //i
    .io_allocateIn_payload_uop_decoded_microcodeEntry                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_microcodeEntry[7:0]          ), //i
    .io_allocateIn_payload_uop_decoded_isSerializing                 (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isSerializing                ), //i
    .io_allocateIn_payload_uop_decoded_isBranchOrJump                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isBranchOrJump               ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_isTaken      (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_isTaken     ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_target       (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_target[31:0]), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted (DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_wasPredicted), //i
    .io_allocateIn_payload_uop_rename_physSrc1_idx                   (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc1_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physSrc1IsFpr                  (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc1IsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_physSrc2_idx                   (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc2_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physSrc2IsFpr                  (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc2IsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_physDest_idx                   (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physDest_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physDestIsFpr                  (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physDestIsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_oldPhysDest_idx                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_oldPhysDest_idx[5:0]          ), //i
    .io_allocateIn_payload_uop_rename_oldPhysDestIsFpr               (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_oldPhysDestIsFpr              ), //i
    .io_allocateIn_payload_uop_rename_allocatesPhysDest              (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_allocatesPhysDest             ), //i
    .io_allocateIn_payload_uop_rename_writesToPhysReg                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_writesToPhysReg               ), //i
    .io_allocateIn_payload_uop_robPtr                                (DispatchPlugin_logic_iqRegs_0_1_payload_uop_robPtr[3:0]                          ), //i
    .io_allocateIn_payload_uop_uniqueId                              (DispatchPlugin_logic_iqRegs_0_1_payload_uop_uniqueId[15:0]                       ), //i
    .io_allocateIn_payload_uop_dispatched                            (DispatchPlugin_logic_iqRegs_0_1_payload_uop_dispatched                           ), //i
    .io_allocateIn_payload_uop_executed                              (DispatchPlugin_logic_iqRegs_0_1_payload_uop_executed                             ), //i
    .io_allocateIn_payload_uop_hasException                          (DispatchPlugin_logic_iqRegs_0_1_payload_uop_hasException                         ), //i
    .io_allocateIn_payload_uop_exceptionCode                         (DispatchPlugin_logic_iqRegs_0_1_payload_uop_exceptionCode[7:0]                   ), //i
    .io_allocateIn_payload_src1InitialReady                          (DispatchPlugin_logic_iqRegs_0_1_payload_src1InitialReady                         ), //i
    .io_allocateIn_payload_src2InitialReady                          (DispatchPlugin_logic_iqRegs_0_1_payload_src2InitialReady                         ), //i
    .io_issueOut_valid                                               (issueQueueComponent_4_io_issueOut_valid                                          ), //o
    .io_issueOut_ready                                               (AluIntEU_AluIntEuPlugin_euInputPort_ready                                        ), //i
    .io_issueOut_payload_robPtr                                      (issueQueueComponent_4_io_issueOut_payload_robPtr[3:0]                            ), //o
    .io_issueOut_payload_physDest_idx                                (issueQueueComponent_4_io_issueOut_payload_physDest_idx[5:0]                      ), //o
    .io_issueOut_payload_physDestIsFpr                               (issueQueueComponent_4_io_issueOut_payload_physDestIsFpr                          ), //o
    .io_issueOut_payload_writesToPhysReg                             (issueQueueComponent_4_io_issueOut_payload_writesToPhysReg                        ), //o
    .io_issueOut_payload_useSrc1                                     (issueQueueComponent_4_io_issueOut_payload_useSrc1                                ), //o
    .io_issueOut_payload_src1Data                                    (issueQueueComponent_4_io_issueOut_payload_src1Data[31:0]                         ), //o
    .io_issueOut_payload_src1Tag                                     (issueQueueComponent_4_io_issueOut_payload_src1Tag[5:0]                           ), //o
    .io_issueOut_payload_src1Ready                                   (issueQueueComponent_4_io_issueOut_payload_src1Ready                              ), //o
    .io_issueOut_payload_src1IsFpr                                   (issueQueueComponent_4_io_issueOut_payload_src1IsFpr                              ), //o
    .io_issueOut_payload_useSrc2                                     (issueQueueComponent_4_io_issueOut_payload_useSrc2                                ), //o
    .io_issueOut_payload_src2Data                                    (issueQueueComponent_4_io_issueOut_payload_src2Data[31:0]                         ), //o
    .io_issueOut_payload_src2Tag                                     (issueQueueComponent_4_io_issueOut_payload_src2Tag[5:0]                           ), //o
    .io_issueOut_payload_src2Ready                                   (issueQueueComponent_4_io_issueOut_payload_src2Ready                              ), //o
    .io_issueOut_payload_src2IsFpr                                   (issueQueueComponent_4_io_issueOut_payload_src2IsFpr                              ), //o
    .io_issueOut_payload_aluCtrl_valid                               (issueQueueComponent_4_io_issueOut_payload_aluCtrl_valid                          ), //o
    .io_issueOut_payload_aluCtrl_isSub                               (issueQueueComponent_4_io_issueOut_payload_aluCtrl_isSub                          ), //o
    .io_issueOut_payload_aluCtrl_isAdd                               (issueQueueComponent_4_io_issueOut_payload_aluCtrl_isAdd                          ), //o
    .io_issueOut_payload_aluCtrl_isSigned                            (issueQueueComponent_4_io_issueOut_payload_aluCtrl_isSigned                       ), //o
    .io_issueOut_payload_aluCtrl_logicOp                             (issueQueueComponent_4_io_issueOut_payload_aluCtrl_logicOp[1:0]                   ), //o
    .io_issueOut_payload_shiftCtrl_valid                             (issueQueueComponent_4_io_issueOut_payload_shiftCtrl_valid                        ), //o
    .io_issueOut_payload_shiftCtrl_isRight                           (issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isRight                      ), //o
    .io_issueOut_payload_shiftCtrl_isArithmetic                      (issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isArithmetic                 ), //o
    .io_issueOut_payload_shiftCtrl_isRotate                          (issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isRotate                     ), //o
    .io_issueOut_payload_shiftCtrl_isDoubleWord                      (issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isDoubleWord                 ), //o
    .io_issueOut_payload_imm                                         (issueQueueComponent_4_io_issueOut_payload_imm[31:0]                              ), //o
    .io_issueOut_payload_immUsage                                    (issueQueueComponent_4_io_issueOut_payload_immUsage[2:0]                          ), //o
    .io_wakeupIn_0_valid                                             (LinkerPlugin_logic_allWakeupFlows_0_valid                                        ), //i
    .io_wakeupIn_0_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_0_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_1_valid                                             (LinkerPlugin_logic_allWakeupFlows_1_valid                                        ), //i
    .io_wakeupIn_1_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_1_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_2_valid                                             (LinkerPlugin_logic_allWakeupFlows_2_valid                                        ), //i
    .io_wakeupIn_2_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_2_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_3_valid                                             (LinkerPlugin_logic_allWakeupFlows_3_valid                                        ), //i
    .io_wakeupIn_3_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_3_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_4_valid                                             (LinkerPlugin_logic_allWakeupFlows_4_valid                                        ), //i
    .io_wakeupIn_4_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_4_payload_physRegIdx[5:0]                      ), //i
    .io_flush                                                        (FetchPipelinePlugin_doHardRedirect_listening                                     ), //i
    .clk                                                             (clk                                                                              ), //i
    .reset                                                           (reset                                                                            )  //i
  );
  IssueQueueComponent_1 issueQueueComponent_5 (
    .io_allocateIn_valid                                             (DispatchPlugin_logic_iqRegs_1_1_valid                                              ), //i
    .io_allocateIn_ready                                             (issueQueueComponent_5_io_allocateIn_ready                                          ), //o
    .io_allocateIn_payload_uop_decoded_pc                            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_pc[31:0]                       ), //i
    .io_allocateIn_payload_uop_decoded_isValid                       (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isValid                        ), //i
    .io_allocateIn_payload_uop_decoded_uopCode                       (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode[4:0]                   ), //i
    .io_allocateIn_payload_uop_decoded_exeUnit                       (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit[3:0]                   ), //i
    .io_allocateIn_payload_uop_decoded_isa                           (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa[1:0]                       ), //i
    .io_allocateIn_payload_uop_decoded_archDest_idx                  (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_idx[4:0]              ), //i
    .io_allocateIn_payload_uop_decoded_archDest_rtype                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype[1:0]            ), //i
    .io_allocateIn_payload_uop_decoded_writeArchDestEn               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_writeArchDestEn                ), //i
    .io_allocateIn_payload_uop_decoded_archSrc1_idx                  (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_idx[4:0]              ), //i
    .io_allocateIn_payload_uop_decoded_archSrc1_rtype                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype[1:0]            ), //i
    .io_allocateIn_payload_uop_decoded_useArchSrc1                   (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_useArchSrc1                    ), //i
    .io_allocateIn_payload_uop_decoded_archSrc2_idx                  (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_idx[4:0]              ), //i
    .io_allocateIn_payload_uop_decoded_archSrc2_rtype                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype[1:0]            ), //i
    .io_allocateIn_payload_uop_decoded_useArchSrc2                   (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_useArchSrc2                    ), //i
    .io_allocateIn_payload_uop_decoded_usePcForAddr                  (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_usePcForAddr                   ), //i
    .io_allocateIn_payload_uop_decoded_imm                           (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_imm[31:0]                      ), //i
    .io_allocateIn_payload_uop_decoded_immUsage                      (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage[2:0]                  ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_valid                 (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_valid                  ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isSub                 (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isSub                  ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isAdd                 (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isAdd                  ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isSigned              (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isSigned               ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_logicOp               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp[1:0]           ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_valid               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_valid                ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isRight             (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isRight              ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic        (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isArithmetic         ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isRotate             ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord        (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isDoubleWord         ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_valid              (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_valid               ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv              (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isDiv               ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned           (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isSigned            ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp           (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isWordOp            ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_size                  (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size[1:0]              ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad          (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isSignedLoad           ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isStore               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isStore                ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked          (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isLoadLinked           ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond           (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isStoreCond            ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_atomicOp              (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_atomicOp[4:0]          ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isFence               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isFence                ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_fenceMode             (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_fenceMode[7:0]         ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp             (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isCacheOp              ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType           (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_cacheOpType[4:0]       ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isPrefetch             ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_condition          (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition[4:0]      ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isJump             (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isJump              ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isLink             (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isLink              ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx        (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_idx[4:0]    ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype      (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype[1:0]  ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect         (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isIndirect          ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_laCfIdx[2:0]        ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_opType                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_opType[3:0]            ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1[1:0]        ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2[1:0]        ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest[1:0]        ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode          (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_roundingMode[2:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest         (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_isIntegerDest          ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt           (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_isSignedCvt            ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1             ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond              (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fcmpCond[4:0]          ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_csrAddr[13:0]          ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isWrite               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isWrite                ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isRead                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isRead                 ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isExchange            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isExchange             ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc          (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_useUimmAsSrc           ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_sysCode               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_sysCode[19:0]          ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn     (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_isExceptionReturn      ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_isTlbOp                ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType             (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_tlbOpType[3:0]         ), //i
    .io_allocateIn_payload_uop_decoded_decodeExceptionCode           (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode[1:0]       ), //i
    .io_allocateIn_payload_uop_decoded_hasDecodeException            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_hasDecodeException             ), //i
    .io_allocateIn_payload_uop_decoded_isMicrocode                   (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isMicrocode                    ), //i
    .io_allocateIn_payload_uop_decoded_microcodeEntry                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_microcodeEntry[7:0]            ), //i
    .io_allocateIn_payload_uop_decoded_isSerializing                 (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isSerializing                  ), //i
    .io_allocateIn_payload_uop_decoded_isBranchOrJump                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isBranchOrJump                 ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_isTaken      (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_isTaken       ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_target       (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_target[31:0]  ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted (DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_wasPredicted  ), //i
    .io_allocateIn_payload_uop_rename_physSrc1_idx                   (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc1_idx[5:0]               ), //i
    .io_allocateIn_payload_uop_rename_physSrc1IsFpr                  (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc1IsFpr                   ), //i
    .io_allocateIn_payload_uop_rename_physSrc2_idx                   (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc2_idx[5:0]               ), //i
    .io_allocateIn_payload_uop_rename_physSrc2IsFpr                  (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc2IsFpr                   ), //i
    .io_allocateIn_payload_uop_rename_physDest_idx                   (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physDest_idx[5:0]               ), //i
    .io_allocateIn_payload_uop_rename_physDestIsFpr                  (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physDestIsFpr                   ), //i
    .io_allocateIn_payload_uop_rename_oldPhysDest_idx                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_oldPhysDest_idx[5:0]            ), //i
    .io_allocateIn_payload_uop_rename_oldPhysDestIsFpr               (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_oldPhysDestIsFpr                ), //i
    .io_allocateIn_payload_uop_rename_allocatesPhysDest              (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_allocatesPhysDest               ), //i
    .io_allocateIn_payload_uop_rename_writesToPhysReg                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_writesToPhysReg                 ), //i
    .io_allocateIn_payload_uop_robPtr                                (DispatchPlugin_logic_iqRegs_1_1_payload_uop_robPtr[3:0]                            ), //i
    .io_allocateIn_payload_uop_uniqueId                              (DispatchPlugin_logic_iqRegs_1_1_payload_uop_uniqueId[15:0]                         ), //i
    .io_allocateIn_payload_uop_dispatched                            (DispatchPlugin_logic_iqRegs_1_1_payload_uop_dispatched                             ), //i
    .io_allocateIn_payload_uop_executed                              (DispatchPlugin_logic_iqRegs_1_1_payload_uop_executed                               ), //i
    .io_allocateIn_payload_uop_hasException                          (DispatchPlugin_logic_iqRegs_1_1_payload_uop_hasException                           ), //i
    .io_allocateIn_payload_uop_exceptionCode                         (DispatchPlugin_logic_iqRegs_1_1_payload_uop_exceptionCode[7:0]                     ), //i
    .io_allocateIn_payload_src1InitialReady                          (DispatchPlugin_logic_iqRegs_1_1_payload_src1InitialReady                           ), //i
    .io_allocateIn_payload_src2InitialReady                          (DispatchPlugin_logic_iqRegs_1_1_payload_src2InitialReady                           ), //i
    .io_issueOut_valid                                               (issueQueueComponent_5_io_issueOut_valid                                            ), //o
    .io_issueOut_ready                                               (MulEU_MulEuPlugin_euInputPort_ready                                                ), //i
    .io_issueOut_payload_uop_decoded_pc                              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_pc[31:0]                     ), //o
    .io_issueOut_payload_uop_decoded_isValid                         (issueQueueComponent_5_io_issueOut_payload_uop_decoded_isValid                      ), //o
    .io_issueOut_payload_uop_decoded_uopCode                         (issueQueueComponent_5_io_issueOut_payload_uop_decoded_uopCode[4:0]                 ), //o
    .io_issueOut_payload_uop_decoded_exeUnit                         (issueQueueComponent_5_io_issueOut_payload_uop_decoded_exeUnit[3:0]                 ), //o
    .io_issueOut_payload_uop_decoded_isa                             (issueQueueComponent_5_io_issueOut_payload_uop_decoded_isa[1:0]                     ), //o
    .io_issueOut_payload_uop_decoded_archDest_idx                    (issueQueueComponent_5_io_issueOut_payload_uop_decoded_archDest_idx[4:0]            ), //o
    .io_issueOut_payload_uop_decoded_archDest_rtype                  (issueQueueComponent_5_io_issueOut_payload_uop_decoded_archDest_rtype[1:0]          ), //o
    .io_issueOut_payload_uop_decoded_writeArchDestEn                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_writeArchDestEn              ), //o
    .io_issueOut_payload_uop_decoded_archSrc1_idx                    (issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc1_idx[4:0]            ), //o
    .io_issueOut_payload_uop_decoded_archSrc1_rtype                  (issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc1_rtype[1:0]          ), //o
    .io_issueOut_payload_uop_decoded_useArchSrc1                     (issueQueueComponent_5_io_issueOut_payload_uop_decoded_useArchSrc1                  ), //o
    .io_issueOut_payload_uop_decoded_archSrc2_idx                    (issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc2_idx[4:0]            ), //o
    .io_issueOut_payload_uop_decoded_archSrc2_rtype                  (issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc2_rtype[1:0]          ), //o
    .io_issueOut_payload_uop_decoded_useArchSrc2                     (issueQueueComponent_5_io_issueOut_payload_uop_decoded_useArchSrc2                  ), //o
    .io_issueOut_payload_uop_decoded_usePcForAddr                    (issueQueueComponent_5_io_issueOut_payload_uop_decoded_usePcForAddr                 ), //o
    .io_issueOut_payload_uop_decoded_imm                             (issueQueueComponent_5_io_issueOut_payload_uop_decoded_imm[31:0]                    ), //o
    .io_issueOut_payload_uop_decoded_immUsage                        (issueQueueComponent_5_io_issueOut_payload_uop_decoded_immUsage[2:0]                ), //o
    .io_issueOut_payload_uop_decoded_aluCtrl_valid                   (issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_valid                ), //o
    .io_issueOut_payload_uop_decoded_aluCtrl_isSub                   (issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isSub                ), //o
    .io_issueOut_payload_uop_decoded_aluCtrl_isAdd                   (issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isAdd                ), //o
    .io_issueOut_payload_uop_decoded_aluCtrl_isSigned                (issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isSigned             ), //o
    .io_issueOut_payload_uop_decoded_aluCtrl_logicOp                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_logicOp[1:0]         ), //o
    .io_issueOut_payload_uop_decoded_shiftCtrl_valid                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_valid              ), //o
    .io_issueOut_payload_uop_decoded_shiftCtrl_isRight               (issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isRight            ), //o
    .io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic          (issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic       ), //o
    .io_issueOut_payload_uop_decoded_shiftCtrl_isRotate              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate           ), //o
    .io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord          (issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord       ), //o
    .io_issueOut_payload_uop_decoded_mulDivCtrl_valid                (issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_valid             ), //o
    .io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv                (issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv             ), //o
    .io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned             (issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned          ), //o
    .io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp             (issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp          ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_size                    (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_size[1:0]            ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad            (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad         ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_isStore                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isStore              ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked            (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked         ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_isStoreCond             (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond          ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_atomicOp                (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_atomicOp[4:0]        ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_isFence                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isFence              ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_fenceMode               (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_fenceMode[7:0]       ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_isCacheOp               (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp            ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_cacheOpType             (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType[4:0]     ), //o
    .io_issueOut_payload_uop_decoded_memCtrl_isPrefetch              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch           ), //o
    .io_issueOut_payload_uop_decoded_branchCtrl_condition            (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_condition[4:0]    ), //o
    .io_issueOut_payload_uop_decoded_branchCtrl_isJump               (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isJump            ), //o
    .io_issueOut_payload_uop_decoded_branchCtrl_isLink               (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isLink            ), //o
    .io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx          (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx[4:0]  ), //o
    .io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype        (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype[1:0]), //o
    .io_issueOut_payload_uop_decoded_branchCtrl_isIndirect           (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect        ), //o
    .io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx[2:0]      ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_opType                  (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_opType[3:0]          ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1[1:0]      ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2[1:0]      ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest[1:0]      ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode            (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode[2:0]    ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest           (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest        ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt             (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt          ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1           ), //o
    .io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond                (issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond[4:0]        ), //o
    .io_issueOut_payload_uop_decoded_csrCtrl_csrAddr                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr[13:0]        ), //o
    .io_issueOut_payload_uop_decoded_csrCtrl_isWrite                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isWrite              ), //o
    .io_issueOut_payload_uop_decoded_csrCtrl_isRead                  (issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isRead               ), //o
    .io_issueOut_payload_uop_decoded_csrCtrl_isExchange              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isExchange           ), //o
    .io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc            (issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc         ), //o
    .io_issueOut_payload_uop_decoded_sysCtrl_sysCode                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_sysCode[19:0]        ), //o
    .io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn       (issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn    ), //o
    .io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp                 (issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp              ), //o
    .io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType               (issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType[3:0]       ), //o
    .io_issueOut_payload_uop_decoded_decodeExceptionCode             (issueQueueComponent_5_io_issueOut_payload_uop_decoded_decodeExceptionCode[1:0]     ), //o
    .io_issueOut_payload_uop_decoded_hasDecodeException              (issueQueueComponent_5_io_issueOut_payload_uop_decoded_hasDecodeException           ), //o
    .io_issueOut_payload_uop_decoded_isMicrocode                     (issueQueueComponent_5_io_issueOut_payload_uop_decoded_isMicrocode                  ), //o
    .io_issueOut_payload_uop_decoded_microcodeEntry                  (issueQueueComponent_5_io_issueOut_payload_uop_decoded_microcodeEntry[7:0]          ), //o
    .io_issueOut_payload_uop_decoded_isSerializing                   (issueQueueComponent_5_io_issueOut_payload_uop_decoded_isSerializing                ), //o
    .io_issueOut_payload_uop_decoded_isBranchOrJump                  (issueQueueComponent_5_io_issueOut_payload_uop_decoded_isBranchOrJump               ), //o
    .io_issueOut_payload_uop_decoded_branchPrediction_isTaken        (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_isTaken     ), //o
    .io_issueOut_payload_uop_decoded_branchPrediction_target         (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_target[31:0]), //o
    .io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted   (issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted), //o
    .io_issueOut_payload_uop_rename_physSrc1_idx                     (issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc1_idx[5:0]             ), //o
    .io_issueOut_payload_uop_rename_physSrc1IsFpr                    (issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc1IsFpr                 ), //o
    .io_issueOut_payload_uop_rename_physSrc2_idx                     (issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc2_idx[5:0]             ), //o
    .io_issueOut_payload_uop_rename_physSrc2IsFpr                    (issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc2IsFpr                 ), //o
    .io_issueOut_payload_uop_rename_physDest_idx                     (issueQueueComponent_5_io_issueOut_payload_uop_rename_physDest_idx[5:0]             ), //o
    .io_issueOut_payload_uop_rename_physDestIsFpr                    (issueQueueComponent_5_io_issueOut_payload_uop_rename_physDestIsFpr                 ), //o
    .io_issueOut_payload_uop_rename_oldPhysDest_idx                  (issueQueueComponent_5_io_issueOut_payload_uop_rename_oldPhysDest_idx[5:0]          ), //o
    .io_issueOut_payload_uop_rename_oldPhysDestIsFpr                 (issueQueueComponent_5_io_issueOut_payload_uop_rename_oldPhysDestIsFpr              ), //o
    .io_issueOut_payload_uop_rename_allocatesPhysDest                (issueQueueComponent_5_io_issueOut_payload_uop_rename_allocatesPhysDest             ), //o
    .io_issueOut_payload_uop_rename_writesToPhysReg                  (issueQueueComponent_5_io_issueOut_payload_uop_rename_writesToPhysReg               ), //o
    .io_issueOut_payload_uop_robPtr                                  (issueQueueComponent_5_io_issueOut_payload_uop_robPtr[3:0]                          ), //o
    .io_issueOut_payload_uop_uniqueId                                (issueQueueComponent_5_io_issueOut_payload_uop_uniqueId[15:0]                       ), //o
    .io_issueOut_payload_uop_dispatched                              (issueQueueComponent_5_io_issueOut_payload_uop_dispatched                           ), //o
    .io_issueOut_payload_uop_executed                                (issueQueueComponent_5_io_issueOut_payload_uop_executed                             ), //o
    .io_issueOut_payload_uop_hasException                            (issueQueueComponent_5_io_issueOut_payload_uop_hasException                         ), //o
    .io_issueOut_payload_uop_exceptionCode                           (issueQueueComponent_5_io_issueOut_payload_uop_exceptionCode[7:0]                   ), //o
    .io_issueOut_payload_robPtr                                      (issueQueueComponent_5_io_issueOut_payload_robPtr[3:0]                              ), //o
    .io_issueOut_payload_physDest_idx                                (issueQueueComponent_5_io_issueOut_payload_physDest_idx[5:0]                        ), //o
    .io_issueOut_payload_physDestIsFpr                               (issueQueueComponent_5_io_issueOut_payload_physDestIsFpr                            ), //o
    .io_issueOut_payload_writesToPhysReg                             (issueQueueComponent_5_io_issueOut_payload_writesToPhysReg                          ), //o
    .io_issueOut_payload_useSrc1                                     (issueQueueComponent_5_io_issueOut_payload_useSrc1                                  ), //o
    .io_issueOut_payload_src1Data                                    (issueQueueComponent_5_io_issueOut_payload_src1Data[31:0]                           ), //o
    .io_issueOut_payload_src1Tag                                     (issueQueueComponent_5_io_issueOut_payload_src1Tag[5:0]                             ), //o
    .io_issueOut_payload_src1Ready                                   (issueQueueComponent_5_io_issueOut_payload_src1Ready                                ), //o
    .io_issueOut_payload_src1IsFpr                                   (issueQueueComponent_5_io_issueOut_payload_src1IsFpr                                ), //o
    .io_issueOut_payload_useSrc2                                     (issueQueueComponent_5_io_issueOut_payload_useSrc2                                  ), //o
    .io_issueOut_payload_src2Data                                    (issueQueueComponent_5_io_issueOut_payload_src2Data[31:0]                           ), //o
    .io_issueOut_payload_src2Tag                                     (issueQueueComponent_5_io_issueOut_payload_src2Tag[5:0]                             ), //o
    .io_issueOut_payload_src2Ready                                   (issueQueueComponent_5_io_issueOut_payload_src2Ready                                ), //o
    .io_issueOut_payload_src2IsFpr                                   (issueQueueComponent_5_io_issueOut_payload_src2IsFpr                                ), //o
    .io_issueOut_payload_mulDivCtrl_valid                            (issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_valid                         ), //o
    .io_issueOut_payload_mulDivCtrl_isDiv                            (issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isDiv                         ), //o
    .io_issueOut_payload_mulDivCtrl_isSigned                         (issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isSigned                      ), //o
    .io_issueOut_payload_mulDivCtrl_isWordOp                         (issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isWordOp                      ), //o
    .io_wakeupIn_0_valid                                             (LinkerPlugin_logic_allWakeupFlows_0_valid                                          ), //i
    .io_wakeupIn_0_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_0_payload_physRegIdx[5:0]                        ), //i
    .io_wakeupIn_1_valid                                             (LinkerPlugin_logic_allWakeupFlows_1_valid                                          ), //i
    .io_wakeupIn_1_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_1_payload_physRegIdx[5:0]                        ), //i
    .io_wakeupIn_2_valid                                             (LinkerPlugin_logic_allWakeupFlows_2_valid                                          ), //i
    .io_wakeupIn_2_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_2_payload_physRegIdx[5:0]                        ), //i
    .io_wakeupIn_3_valid                                             (LinkerPlugin_logic_allWakeupFlows_3_valid                                          ), //i
    .io_wakeupIn_3_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_3_payload_physRegIdx[5:0]                        ), //i
    .io_wakeupIn_4_valid                                             (LinkerPlugin_logic_allWakeupFlows_4_valid                                          ), //i
    .io_wakeupIn_4_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_4_payload_physRegIdx[5:0]                        ), //i
    .io_flush                                                        (FetchPipelinePlugin_doHardRedirect_listening                                       ), //i
    .clk                                                             (clk                                                                                ), //i
    .reset                                                           (reset                                                                              )  //i
  );
  IssueQueueComponent_2 issueQueueComponent_6 (
    .io_allocateIn_valid                                             (DispatchPlugin_logic_iqRegs_2_1_valid                                            ), //i
    .io_allocateIn_ready                                             (issueQueueComponent_6_io_allocateIn_ready                                        ), //o
    .io_allocateIn_payload_uop_decoded_pc                            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_pc[31:0]                     ), //i
    .io_allocateIn_payload_uop_decoded_isValid                       (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isValid                      ), //i
    .io_allocateIn_payload_uop_decoded_uopCode                       (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode[4:0]                 ), //i
    .io_allocateIn_payload_uop_decoded_exeUnit                       (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit[3:0]                 ), //i
    .io_allocateIn_payload_uop_decoded_isa                           (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa[1:0]                     ), //i
    .io_allocateIn_payload_uop_decoded_archDest_idx                  (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archDest_rtype                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_writeArchDestEn               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_writeArchDestEn              ), //i
    .io_allocateIn_payload_uop_decoded_archSrc1_idx                  (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archSrc1_rtype                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_useArchSrc1                   (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_useArchSrc1                  ), //i
    .io_allocateIn_payload_uop_decoded_archSrc2_idx                  (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archSrc2_rtype                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_useArchSrc2                   (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_useArchSrc2                  ), //i
    .io_allocateIn_payload_uop_decoded_usePcForAddr                  (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_usePcForAddr                 ), //i
    .io_allocateIn_payload_uop_decoded_imm                           (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_imm[31:0]                    ), //i
    .io_allocateIn_payload_uop_decoded_immUsage                      (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage[2:0]                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_valid                 (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_valid                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isSub                 (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isSub                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isAdd                 (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isAdd                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isSigned              (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isSigned             ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_logicOp               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp[1:0]         ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_valid               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_valid              ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isRight             (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isRight            ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic        (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isArithmetic       ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isRotate           ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord        (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isDoubleWord       ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_valid              (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_valid             ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv              (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isDiv             ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned           (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isSigned          ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp           (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isWordOp          ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_size                  (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size[1:0]            ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad          (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isSignedLoad         ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isStore               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isStore              ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked          (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isLoadLinked         ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond           (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isStoreCond          ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_atomicOp              (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_atomicOp[4:0]        ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isFence               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isFence              ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_fenceMode             (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_fenceMode[7:0]       ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp             (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isCacheOp            ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType           (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_cacheOpType[4:0]     ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isPrefetch           ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_condition          (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition[4:0]    ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isJump             (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isJump            ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isLink             (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isLink            ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx        (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_idx[4:0]  ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype      (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype[1:0]), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect         (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isIndirect        ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_laCfIdx[2:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_opType                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_opType[3:0]          ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode          (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_roundingMode[2:0]    ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest         (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_isIntegerDest        ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt           (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_isSignedCvt          ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1           ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond              (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fcmpCond[4:0]        ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_csrAddr[13:0]        ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isWrite               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isWrite              ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isRead                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isRead               ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isExchange            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isExchange           ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc          (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_useUimmAsSrc         ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_sysCode               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_sysCode[19:0]        ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn     (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_isExceptionReturn    ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_isTlbOp              ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType             (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_tlbOpType[3:0]       ), //i
    .io_allocateIn_payload_uop_decoded_decodeExceptionCode           (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode[1:0]     ), //i
    .io_allocateIn_payload_uop_decoded_hasDecodeException            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_hasDecodeException           ), //i
    .io_allocateIn_payload_uop_decoded_isMicrocode                   (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isMicrocode                  ), //i
    .io_allocateIn_payload_uop_decoded_microcodeEntry                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_microcodeEntry[7:0]          ), //i
    .io_allocateIn_payload_uop_decoded_isSerializing                 (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isSerializing                ), //i
    .io_allocateIn_payload_uop_decoded_isBranchOrJump                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isBranchOrJump               ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_isTaken      (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_isTaken     ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_target       (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_target[31:0]), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted (DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_wasPredicted), //i
    .io_allocateIn_payload_uop_rename_physSrc1_idx                   (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc1_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physSrc1IsFpr                  (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc1IsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_physSrc2_idx                   (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc2_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physSrc2IsFpr                  (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc2IsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_physDest_idx                   (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physDest_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physDestIsFpr                  (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physDestIsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_oldPhysDest_idx                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_oldPhysDest_idx[5:0]          ), //i
    .io_allocateIn_payload_uop_rename_oldPhysDestIsFpr               (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_oldPhysDestIsFpr              ), //i
    .io_allocateIn_payload_uop_rename_allocatesPhysDest              (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_allocatesPhysDest             ), //i
    .io_allocateIn_payload_uop_rename_writesToPhysReg                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_writesToPhysReg               ), //i
    .io_allocateIn_payload_uop_robPtr                                (DispatchPlugin_logic_iqRegs_2_1_payload_uop_robPtr[3:0]                          ), //i
    .io_allocateIn_payload_uop_uniqueId                              (DispatchPlugin_logic_iqRegs_2_1_payload_uop_uniqueId[15:0]                       ), //i
    .io_allocateIn_payload_uop_dispatched                            (DispatchPlugin_logic_iqRegs_2_1_payload_uop_dispatched                           ), //i
    .io_allocateIn_payload_uop_executed                              (DispatchPlugin_logic_iqRegs_2_1_payload_uop_executed                             ), //i
    .io_allocateIn_payload_uop_hasException                          (DispatchPlugin_logic_iqRegs_2_1_payload_uop_hasException                         ), //i
    .io_allocateIn_payload_uop_exceptionCode                         (DispatchPlugin_logic_iqRegs_2_1_payload_uop_exceptionCode[7:0]                   ), //i
    .io_allocateIn_payload_src1InitialReady                          (DispatchPlugin_logic_iqRegs_2_1_payload_src1InitialReady                         ), //i
    .io_allocateIn_payload_src2InitialReady                          (DispatchPlugin_logic_iqRegs_2_1_payload_src2InitialReady                         ), //i
    .io_issueOut_valid                                               (issueQueueComponent_6_io_issueOut_valid                                          ), //o
    .io_issueOut_ready                                               (BranchEU_BranchEuPlugin_euInputPort_ready                                        ), //i
    .io_issueOut_payload_robPtr                                      (issueQueueComponent_6_io_issueOut_payload_robPtr[3:0]                            ), //o
    .io_issueOut_payload_physDest_idx                                (issueQueueComponent_6_io_issueOut_payload_physDest_idx[5:0]                      ), //o
    .io_issueOut_payload_physDestIsFpr                               (issueQueueComponent_6_io_issueOut_payload_physDestIsFpr                          ), //o
    .io_issueOut_payload_writesToPhysReg                             (issueQueueComponent_6_io_issueOut_payload_writesToPhysReg                        ), //o
    .io_issueOut_payload_useSrc1                                     (issueQueueComponent_6_io_issueOut_payload_useSrc1                                ), //o
    .io_issueOut_payload_src1Data                                    (issueQueueComponent_6_io_issueOut_payload_src1Data[31:0]                         ), //o
    .io_issueOut_payload_src1Tag                                     (issueQueueComponent_6_io_issueOut_payload_src1Tag[5:0]                           ), //o
    .io_issueOut_payload_src1Ready                                   (issueQueueComponent_6_io_issueOut_payload_src1Ready                              ), //o
    .io_issueOut_payload_src1IsFpr                                   (issueQueueComponent_6_io_issueOut_payload_src1IsFpr                              ), //o
    .io_issueOut_payload_useSrc2                                     (issueQueueComponent_6_io_issueOut_payload_useSrc2                                ), //o
    .io_issueOut_payload_src2Data                                    (issueQueueComponent_6_io_issueOut_payload_src2Data[31:0]                         ), //o
    .io_issueOut_payload_src2Tag                                     (issueQueueComponent_6_io_issueOut_payload_src2Tag[5:0]                           ), //o
    .io_issueOut_payload_src2Ready                                   (issueQueueComponent_6_io_issueOut_payload_src2Ready                              ), //o
    .io_issueOut_payload_src2IsFpr                                   (issueQueueComponent_6_io_issueOut_payload_src2IsFpr                              ), //o
    .io_issueOut_payload_branchCtrl_condition                        (issueQueueComponent_6_io_issueOut_payload_branchCtrl_condition[4:0]              ), //o
    .io_issueOut_payload_branchCtrl_isJump                           (issueQueueComponent_6_io_issueOut_payload_branchCtrl_isJump                      ), //o
    .io_issueOut_payload_branchCtrl_isLink                           (issueQueueComponent_6_io_issueOut_payload_branchCtrl_isLink                      ), //o
    .io_issueOut_payload_branchCtrl_linkReg_idx                      (issueQueueComponent_6_io_issueOut_payload_branchCtrl_linkReg_idx[4:0]            ), //o
    .io_issueOut_payload_branchCtrl_linkReg_rtype                    (issueQueueComponent_6_io_issueOut_payload_branchCtrl_linkReg_rtype[1:0]          ), //o
    .io_issueOut_payload_branchCtrl_isIndirect                       (issueQueueComponent_6_io_issueOut_payload_branchCtrl_isIndirect                  ), //o
    .io_issueOut_payload_branchCtrl_laCfIdx                          (issueQueueComponent_6_io_issueOut_payload_branchCtrl_laCfIdx[2:0]                ), //o
    .io_issueOut_payload_imm                                         (issueQueueComponent_6_io_issueOut_payload_imm[31:0]                              ), //o
    .io_issueOut_payload_pc                                          (issueQueueComponent_6_io_issueOut_payload_pc[31:0]                               ), //o
    .io_issueOut_payload_branchPrediction_isTaken                    (issueQueueComponent_6_io_issueOut_payload_branchPrediction_isTaken               ), //o
    .io_issueOut_payload_branchPrediction_target                     (issueQueueComponent_6_io_issueOut_payload_branchPrediction_target[31:0]          ), //o
    .io_issueOut_payload_branchPrediction_wasPredicted               (issueQueueComponent_6_io_issueOut_payload_branchPrediction_wasPredicted          ), //o
    .io_wakeupIn_0_valid                                             (LinkerPlugin_logic_allWakeupFlows_0_valid                                        ), //i
    .io_wakeupIn_0_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_0_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_1_valid                                             (LinkerPlugin_logic_allWakeupFlows_1_valid                                        ), //i
    .io_wakeupIn_1_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_1_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_2_valid                                             (LinkerPlugin_logic_allWakeupFlows_2_valid                                        ), //i
    .io_wakeupIn_2_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_2_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_3_valid                                             (LinkerPlugin_logic_allWakeupFlows_3_valid                                        ), //i
    .io_wakeupIn_3_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_3_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_4_valid                                             (LinkerPlugin_logic_allWakeupFlows_4_valid                                        ), //i
    .io_wakeupIn_4_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_4_payload_physRegIdx[5:0]                      ), //i
    .io_flush                                                        (FetchPipelinePlugin_doHardRedirect_listening                                     ), //i
    .clk                                                             (clk                                                                              ), //i
    .reset                                                           (reset                                                                            )  //i
  );
  IssueQueueComponent_3 issueQueueComponent_7 (
    .io_allocateIn_valid                                             (DispatchPlugin_logic_iqRegs_3_1_valid                                            ), //i
    .io_allocateIn_ready                                             (issueQueueComponent_7_io_allocateIn_ready                                        ), //o
    .io_allocateIn_payload_uop_decoded_pc                            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_pc[31:0]                     ), //i
    .io_allocateIn_payload_uop_decoded_isValid                       (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isValid                      ), //i
    .io_allocateIn_payload_uop_decoded_uopCode                       (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode[4:0]                 ), //i
    .io_allocateIn_payload_uop_decoded_exeUnit                       (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit[3:0]                 ), //i
    .io_allocateIn_payload_uop_decoded_isa                           (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa[1:0]                     ), //i
    .io_allocateIn_payload_uop_decoded_archDest_idx                  (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archDest_rtype                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_writeArchDestEn               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_writeArchDestEn              ), //i
    .io_allocateIn_payload_uop_decoded_archSrc1_idx                  (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archSrc1_rtype                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_useArchSrc1                   (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_useArchSrc1                  ), //i
    .io_allocateIn_payload_uop_decoded_archSrc2_idx                  (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_idx[4:0]            ), //i
    .io_allocateIn_payload_uop_decoded_archSrc2_rtype                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype[1:0]          ), //i
    .io_allocateIn_payload_uop_decoded_useArchSrc2                   (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_useArchSrc2                  ), //i
    .io_allocateIn_payload_uop_decoded_usePcForAddr                  (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_usePcForAddr                 ), //i
    .io_allocateIn_payload_uop_decoded_imm                           (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_imm[31:0]                    ), //i
    .io_allocateIn_payload_uop_decoded_immUsage                      (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage[2:0]                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_valid                 (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_valid                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isSub                 (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isSub                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isAdd                 (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isAdd                ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_isSigned              (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isSigned             ), //i
    .io_allocateIn_payload_uop_decoded_aluCtrl_logicOp               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp[1:0]         ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_valid               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_valid              ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isRight             (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isRight            ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic        (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isArithmetic       ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isRotate           ), //i
    .io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord        (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isDoubleWord       ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_valid              (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_valid             ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv              (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isDiv             ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned           (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isSigned          ), //i
    .io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp           (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isWordOp          ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_size                  (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size[1:0]            ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad          (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isSignedLoad         ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isStore               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isStore              ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked          (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isLoadLinked         ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond           (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isStoreCond          ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_atomicOp              (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_atomicOp[4:0]        ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isFence               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isFence              ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_fenceMode             (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_fenceMode[7:0]       ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp             (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isCacheOp            ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType           (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_cacheOpType[4:0]     ), //i
    .io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isPrefetch           ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_condition          (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition[4:0]    ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isJump             (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isJump            ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isLink             (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isLink            ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx        (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_idx[4:0]  ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype      (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype[1:0]), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect         (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isIndirect        ), //i
    .io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_laCfIdx[2:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_opType                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_opType[3:0]          ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest[1:0]      ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode          (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_roundingMode[2:0]    ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest         (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_isIntegerDest        ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt           (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_isSignedCvt          ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1           ), //i
    .io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond              (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fcmpCond[4:0]        ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_csrAddr[13:0]        ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isWrite               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isWrite              ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isRead                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isRead               ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_isExchange            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isExchange           ), //i
    .io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc          (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_useUimmAsSrc         ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_sysCode               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_sysCode[19:0]        ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn     (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_isExceptionReturn    ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_isTlbOp              ), //i
    .io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType             (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_tlbOpType[3:0]       ), //i
    .io_allocateIn_payload_uop_decoded_decodeExceptionCode           (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode[1:0]     ), //i
    .io_allocateIn_payload_uop_decoded_hasDecodeException            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_hasDecodeException           ), //i
    .io_allocateIn_payload_uop_decoded_isMicrocode                   (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isMicrocode                  ), //i
    .io_allocateIn_payload_uop_decoded_microcodeEntry                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_microcodeEntry[7:0]          ), //i
    .io_allocateIn_payload_uop_decoded_isSerializing                 (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isSerializing                ), //i
    .io_allocateIn_payload_uop_decoded_isBranchOrJump                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isBranchOrJump               ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_isTaken      (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_isTaken     ), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_target       (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_target[31:0]), //i
    .io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted (DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_wasPredicted), //i
    .io_allocateIn_payload_uop_rename_physSrc1_idx                   (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc1_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physSrc1IsFpr                  (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc1IsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_physSrc2_idx                   (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc2_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physSrc2IsFpr                  (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc2IsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_physDest_idx                   (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physDest_idx[5:0]             ), //i
    .io_allocateIn_payload_uop_rename_physDestIsFpr                  (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physDestIsFpr                 ), //i
    .io_allocateIn_payload_uop_rename_oldPhysDest_idx                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_oldPhysDest_idx[5:0]          ), //i
    .io_allocateIn_payload_uop_rename_oldPhysDestIsFpr               (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_oldPhysDestIsFpr              ), //i
    .io_allocateIn_payload_uop_rename_allocatesPhysDest              (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_allocatesPhysDest             ), //i
    .io_allocateIn_payload_uop_rename_writesToPhysReg                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_writesToPhysReg               ), //i
    .io_allocateIn_payload_uop_robPtr                                (DispatchPlugin_logic_iqRegs_3_1_payload_uop_robPtr[3:0]                          ), //i
    .io_allocateIn_payload_uop_uniqueId                              (DispatchPlugin_logic_iqRegs_3_1_payload_uop_uniqueId[15:0]                       ), //i
    .io_allocateIn_payload_uop_dispatched                            (DispatchPlugin_logic_iqRegs_3_1_payload_uop_dispatched                           ), //i
    .io_allocateIn_payload_uop_executed                              (DispatchPlugin_logic_iqRegs_3_1_payload_uop_executed                             ), //i
    .io_allocateIn_payload_uop_hasException                          (DispatchPlugin_logic_iqRegs_3_1_payload_uop_hasException                         ), //i
    .io_allocateIn_payload_uop_exceptionCode                         (DispatchPlugin_logic_iqRegs_3_1_payload_uop_exceptionCode[7:0]                   ), //i
    .io_allocateIn_payload_src1InitialReady                          (DispatchPlugin_logic_iqRegs_3_1_payload_src1InitialReady                         ), //i
    .io_allocateIn_payload_src2InitialReady                          (DispatchPlugin_logic_iqRegs_3_1_payload_src2InitialReady                         ), //i
    .io_issueOut_valid                                               (issueQueueComponent_7_io_issueOut_valid                                          ), //o
    .io_issueOut_ready                                               (LsuEU_LsuEuPlugin_euInputPort_ready                                              ), //i
    .io_issueOut_payload_robPtr                                      (issueQueueComponent_7_io_issueOut_payload_robPtr[3:0]                            ), //o
    .io_issueOut_payload_physDest_idx                                (issueQueueComponent_7_io_issueOut_payload_physDest_idx[5:0]                      ), //o
    .io_issueOut_payload_physDestIsFpr                               (issueQueueComponent_7_io_issueOut_payload_physDestIsFpr                          ), //o
    .io_issueOut_payload_writesToPhysReg                             (issueQueueComponent_7_io_issueOut_payload_writesToPhysReg                        ), //o
    .io_issueOut_payload_useSrc1                                     (issueQueueComponent_7_io_issueOut_payload_useSrc1                                ), //o
    .io_issueOut_payload_src1Data                                    (issueQueueComponent_7_io_issueOut_payload_src1Data[31:0]                         ), //o
    .io_issueOut_payload_src1Tag                                     (issueQueueComponent_7_io_issueOut_payload_src1Tag[5:0]                           ), //o
    .io_issueOut_payload_src1Ready                                   (issueQueueComponent_7_io_issueOut_payload_src1Ready                              ), //o
    .io_issueOut_payload_src1IsFpr                                   (issueQueueComponent_7_io_issueOut_payload_src1IsFpr                              ), //o
    .io_issueOut_payload_useSrc2                                     (issueQueueComponent_7_io_issueOut_payload_useSrc2                                ), //o
    .io_issueOut_payload_src2Data                                    (issueQueueComponent_7_io_issueOut_payload_src2Data[31:0]                         ), //o
    .io_issueOut_payload_src2Tag                                     (issueQueueComponent_7_io_issueOut_payload_src2Tag[5:0]                           ), //o
    .io_issueOut_payload_src2Ready                                   (issueQueueComponent_7_io_issueOut_payload_src2Ready                              ), //o
    .io_issueOut_payload_src2IsFpr                                   (issueQueueComponent_7_io_issueOut_payload_src2IsFpr                              ), //o
    .io_issueOut_payload_memCtrl_size                                (issueQueueComponent_7_io_issueOut_payload_memCtrl_size[1:0]                      ), //o
    .io_issueOut_payload_memCtrl_isSignedLoad                        (issueQueueComponent_7_io_issueOut_payload_memCtrl_isSignedLoad                   ), //o
    .io_issueOut_payload_memCtrl_isStore                             (issueQueueComponent_7_io_issueOut_payload_memCtrl_isStore                        ), //o
    .io_issueOut_payload_memCtrl_isLoadLinked                        (issueQueueComponent_7_io_issueOut_payload_memCtrl_isLoadLinked                   ), //o
    .io_issueOut_payload_memCtrl_isStoreCond                         (issueQueueComponent_7_io_issueOut_payload_memCtrl_isStoreCond                    ), //o
    .io_issueOut_payload_memCtrl_atomicOp                            (issueQueueComponent_7_io_issueOut_payload_memCtrl_atomicOp[4:0]                  ), //o
    .io_issueOut_payload_memCtrl_isFence                             (issueQueueComponent_7_io_issueOut_payload_memCtrl_isFence                        ), //o
    .io_issueOut_payload_memCtrl_fenceMode                           (issueQueueComponent_7_io_issueOut_payload_memCtrl_fenceMode[7:0]                 ), //o
    .io_issueOut_payload_memCtrl_isCacheOp                           (issueQueueComponent_7_io_issueOut_payload_memCtrl_isCacheOp                      ), //o
    .io_issueOut_payload_memCtrl_cacheOpType                         (issueQueueComponent_7_io_issueOut_payload_memCtrl_cacheOpType[4:0]               ), //o
    .io_issueOut_payload_memCtrl_isPrefetch                          (issueQueueComponent_7_io_issueOut_payload_memCtrl_isPrefetch                     ), //o
    .io_issueOut_payload_imm                                         (issueQueueComponent_7_io_issueOut_payload_imm[31:0]                              ), //o
    .io_issueOut_payload_usePc                                       (issueQueueComponent_7_io_issueOut_payload_usePc                                  ), //o
    .io_issueOut_payload_pcData                                      (issueQueueComponent_7_io_issueOut_payload_pcData[31:0]                           ), //o
    .io_wakeupIn_0_valid                                             (LinkerPlugin_logic_allWakeupFlows_0_valid                                        ), //i
    .io_wakeupIn_0_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_0_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_1_valid                                             (LinkerPlugin_logic_allWakeupFlows_1_valid                                        ), //i
    .io_wakeupIn_1_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_1_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_2_valid                                             (LinkerPlugin_logic_allWakeupFlows_2_valid                                        ), //i
    .io_wakeupIn_2_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_2_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_3_valid                                             (LinkerPlugin_logic_allWakeupFlows_3_valid                                        ), //i
    .io_wakeupIn_3_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_3_payload_physRegIdx[5:0]                      ), //i
    .io_wakeupIn_4_valid                                             (LinkerPlugin_logic_allWakeupFlows_4_valid                                        ), //i
    .io_wakeupIn_4_payload_physRegIdx                                (LinkerPlugin_logic_allWakeupFlows_4_payload_physRegIdx[5:0]                      ), //i
    .io_flush                                                        (FetchPipelinePlugin_doHardRedirect_listening                                     ), //i
    .clk                                                             (clk                                                                              ), //i
    .reset                                                           (reset                                                                            )  //i
  );
  OneShot oneShot_20 (
    .io_triggerIn (oneShot_20_io_triggerIn), //i
    .io_pulseOut  (oneShot_20_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  FrequencyDivider DebugDisplayPlugin_logic_displayArea_divider (
    .io_tick (DebugDisplayPlugin_logic_displayArea_divider_io_tick), //o
    .clk     (clk                                                 ), //i
    .reset   (reset                                               )  //i
  );
  OneShot oneShot_21 (
    .io_triggerIn (oneShot_21_io_triggerIn), //i
    .io_pulseOut  (oneShot_21_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  mult_gen_0 multiplierBlackbox (
    .CLK (clk                       ), //i
    .A   (multiplierBlackbox_A[31:0]), //i
    .B   (multiplierBlackbox_B[31:0]), //i
    .P   (multiplierBlackbox_P[63:0])  //o
  );
  OneShot oneShot_22 (
    .io_triggerIn (oneShot_22_io_triggerIn), //i
    .io_pulseOut  (oneShot_22_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  OneShot oneShot_23 (
    .io_triggerIn (oneShot_23_io_triggerIn), //i
    .io_pulseOut  (oneShot_23_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  StreamDemux streamDemux_1 (
    .io_select                           (streamDemux_1_io_select                                     ), //i
    .io_input_valid                      (LsuEU_LsuEuPlugin_hw_aguPort_output_valid                   ), //i
    .io_input_ready                      (streamDemux_1_io_input_ready                                ), //o
    .io_input_payload_qPtr               (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr[2:0]       ), //i
    .io_input_payload_address            (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address[31:0]   ), //i
    .io_input_payload_alignException     (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException  ), //i
    .io_input_payload_accessSize         (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize[1:0] ), //i
    .io_input_payload_storeMask          (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask[3:0]  ), //i
    .io_input_payload_basePhysReg        (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_basePhysReg[5:0]), //i
    .io_input_payload_immediate          (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate[31:0] ), //i
    .io_input_payload_usePc              (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc           ), //i
    .io_input_payload_pc                 (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc[31:0]        ), //i
    .io_input_payload_robPtr             (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr[3:0]     ), //i
    .io_input_payload_isLoad             (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad          ), //i
    .io_input_payload_isStore            (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isStore         ), //i
    .io_input_payload_physDst            (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst[5:0]    ), //i
    .io_input_payload_storeData          (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData[31:0] ), //i
    .io_input_payload_isFlush            (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush         ), //i
    .io_input_payload_isIO               (LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO            ), //i
    .io_outputs_0_valid                  (streamDemux_1_io_outputs_0_valid                            ), //o
    .io_outputs_0_ready                  (io_outputs_0_combStage_ready                                ), //i
    .io_outputs_0_payload_qPtr           (streamDemux_1_io_outputs_0_payload_qPtr[2:0]                ), //o
    .io_outputs_0_payload_address        (streamDemux_1_io_outputs_0_payload_address[31:0]            ), //o
    .io_outputs_0_payload_alignException (streamDemux_1_io_outputs_0_payload_alignException           ), //o
    .io_outputs_0_payload_accessSize     (streamDemux_1_io_outputs_0_payload_accessSize[1:0]          ), //o
    .io_outputs_0_payload_storeMask      (streamDemux_1_io_outputs_0_payload_storeMask[3:0]           ), //o
    .io_outputs_0_payload_basePhysReg    (streamDemux_1_io_outputs_0_payload_basePhysReg[5:0]         ), //o
    .io_outputs_0_payload_immediate      (streamDemux_1_io_outputs_0_payload_immediate[31:0]          ), //o
    .io_outputs_0_payload_usePc          (streamDemux_1_io_outputs_0_payload_usePc                    ), //o
    .io_outputs_0_payload_pc             (streamDemux_1_io_outputs_0_payload_pc[31:0]                 ), //o
    .io_outputs_0_payload_robPtr         (streamDemux_1_io_outputs_0_payload_robPtr[3:0]              ), //o
    .io_outputs_0_payload_isLoad         (streamDemux_1_io_outputs_0_payload_isLoad                   ), //o
    .io_outputs_0_payload_isStore        (streamDemux_1_io_outputs_0_payload_isStore                  ), //o
    .io_outputs_0_payload_physDst        (streamDemux_1_io_outputs_0_payload_physDst[5:0]             ), //o
    .io_outputs_0_payload_storeData      (streamDemux_1_io_outputs_0_payload_storeData[31:0]          ), //o
    .io_outputs_0_payload_isFlush        (streamDemux_1_io_outputs_0_payload_isFlush                  ), //o
    .io_outputs_0_payload_isIO           (streamDemux_1_io_outputs_0_payload_isIO                     ), //o
    .io_outputs_1_valid                  (streamDemux_1_io_outputs_1_valid                            ), //o
    .io_outputs_1_ready                  (io_outputs_1_combStage_ready                                ), //i
    .io_outputs_1_payload_qPtr           (streamDemux_1_io_outputs_1_payload_qPtr[2:0]                ), //o
    .io_outputs_1_payload_address        (streamDemux_1_io_outputs_1_payload_address[31:0]            ), //o
    .io_outputs_1_payload_alignException (streamDemux_1_io_outputs_1_payload_alignException           ), //o
    .io_outputs_1_payload_accessSize     (streamDemux_1_io_outputs_1_payload_accessSize[1:0]          ), //o
    .io_outputs_1_payload_storeMask      (streamDemux_1_io_outputs_1_payload_storeMask[3:0]           ), //o
    .io_outputs_1_payload_basePhysReg    (streamDemux_1_io_outputs_1_payload_basePhysReg[5:0]         ), //o
    .io_outputs_1_payload_immediate      (streamDemux_1_io_outputs_1_payload_immediate[31:0]          ), //o
    .io_outputs_1_payload_usePc          (streamDemux_1_io_outputs_1_payload_usePc                    ), //o
    .io_outputs_1_payload_pc             (streamDemux_1_io_outputs_1_payload_pc[31:0]                 ), //o
    .io_outputs_1_payload_robPtr         (streamDemux_1_io_outputs_1_payload_robPtr[3:0]              ), //o
    .io_outputs_1_payload_isLoad         (streamDemux_1_io_outputs_1_payload_isLoad                   ), //o
    .io_outputs_1_payload_isStore        (streamDemux_1_io_outputs_1_payload_isStore                  ), //o
    .io_outputs_1_payload_physDst        (streamDemux_1_io_outputs_1_payload_physDst[5:0]             ), //o
    .io_outputs_1_payload_storeData      (streamDemux_1_io_outputs_1_payload_storeData[31:0]          ), //o
    .io_outputs_1_payload_isFlush        (streamDemux_1_io_outputs_1_payload_isFlush                  ), //o
    .io_outputs_1_payload_isIO           (streamDemux_1_io_outputs_1_payload_isIO                     )  //o
  );
  OneShot oneShot_24 (
    .io_triggerIn (oneShot_24_io_triggerIn), //i
    .io_pulseOut  (oneShot_24_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  StreamArbiter_7 streamArbiter_9 (
    .io_inputs_0_valid                      (LsuEU_LsuEuPlugin_hw_lqPushPort_valid                          ), //i
    .io_inputs_0_ready                      (streamArbiter_9_io_inputs_0_ready                              ), //o
    .io_inputs_0_payload_robPtr             (LsuEU_LsuEuPlugin_hw_lqPushPort_payload_robPtr[3:0]            ), //i
    .io_inputs_0_payload_pdest              (LsuEU_LsuEuPlugin_hw_lqPushPort_payload_pdest[5:0]             ), //i
    .io_inputs_0_payload_address            (LsuEU_LsuEuPlugin_hw_lqPushPort_payload_address[31:0]          ), //i
    .io_inputs_0_payload_isIO               (LsuEU_LsuEuPlugin_hw_lqPushPort_payload_isIO                   ), //i
    .io_inputs_0_payload_size               (LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size[1:0]              ), //i
    .io_inputs_0_payload_hasEarlyException  (LsuEU_LsuEuPlugin_hw_lqPushPort_payload_hasEarlyException      ), //i
    .io_inputs_0_payload_earlyExceptionCode (LsuEU_LsuEuPlugin_hw_lqPushPort_payload_earlyExceptionCode[7:0]), //i
    .io_output_valid                        (streamArbiter_9_io_output_valid                                ), //o
    .io_output_ready                        (LoadQueuePlugin_logic_pushCmd_ready                            ), //i
    .io_output_payload_robPtr               (streamArbiter_9_io_output_payload_robPtr[3:0]                  ), //o
    .io_output_payload_pdest                (streamArbiter_9_io_output_payload_pdest[5:0]                   ), //o
    .io_output_payload_address              (streamArbiter_9_io_output_payload_address[31:0]                ), //o
    .io_output_payload_isIO                 (streamArbiter_9_io_output_payload_isIO                         ), //o
    .io_output_payload_size                 (streamArbiter_9_io_output_payload_size[1:0]                    ), //o
    .io_output_payload_hasEarlyException    (streamArbiter_9_io_output_payload_hasEarlyException            ), //o
    .io_output_payload_earlyExceptionCode   (streamArbiter_9_io_output_payload_earlyExceptionCode[7:0]      ), //o
    .io_chosenOH                            (streamArbiter_9_io_chosenOH                                    ), //o
    .clk                                    (clk                                                            ), //i
    .reset                                  (reset                                                          )  //i
  );
  OneShot oneShot_25 (
    .io_triggerIn (oneShot_25_io_triggerIn), //i
    .io_pulseOut  (oneShot_25_io_pulseOut ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  SmartDispatcher FetchPipelinePlugin_logic_dispatcher (
    .io_fetchGroupIn_valid                                 (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_valid                                    ), //i
    .io_fetchGroupIn_ready                                 (FetchPipelinePlugin_logic_dispatcher_io_fetchGroupIn_ready                                          ), //o
    .io_fetchGroupIn_payload_pc                            (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_pc[31:0]                         ), //i
    .io_fetchGroupIn_payload_instructions_0                (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_0[31:0]             ), //i
    .io_fetchGroupIn_payload_instructions_1                (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_1[31:0]             ), //i
    .io_fetchGroupIn_payload_instructions_2                (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_2[31:0]             ), //i
    .io_fetchGroupIn_payload_instructions_3                (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_3[31:0]             ), //i
    .io_fetchGroupIn_payload_predecodeInfos_0_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isBranch        ), //i
    .io_fetchGroupIn_payload_predecodeInfos_0_isJump       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isJump          ), //i
    .io_fetchGroupIn_payload_predecodeInfos_0_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isDirectJump    ), //i
    .io_fetchGroupIn_payload_predecodeInfos_0_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_jumpOffset[31:0]), //i
    .io_fetchGroupIn_payload_predecodeInfos_0_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isIdle          ), //i
    .io_fetchGroupIn_payload_predecodeInfos_1_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isBranch        ), //i
    .io_fetchGroupIn_payload_predecodeInfos_1_isJump       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isJump          ), //i
    .io_fetchGroupIn_payload_predecodeInfos_1_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isDirectJump    ), //i
    .io_fetchGroupIn_payload_predecodeInfos_1_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_jumpOffset[31:0]), //i
    .io_fetchGroupIn_payload_predecodeInfos_1_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isIdle          ), //i
    .io_fetchGroupIn_payload_predecodeInfos_2_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isBranch        ), //i
    .io_fetchGroupIn_payload_predecodeInfos_2_isJump       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isJump          ), //i
    .io_fetchGroupIn_payload_predecodeInfos_2_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isDirectJump    ), //i
    .io_fetchGroupIn_payload_predecodeInfos_2_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_jumpOffset[31:0]), //i
    .io_fetchGroupIn_payload_predecodeInfos_2_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isIdle          ), //i
    .io_fetchGroupIn_payload_predecodeInfos_3_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isBranch        ), //i
    .io_fetchGroupIn_payload_predecodeInfos_3_isJump       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isJump          ), //i
    .io_fetchGroupIn_payload_predecodeInfos_3_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isDirectJump    ), //i
    .io_fetchGroupIn_payload_predecodeInfos_3_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_jumpOffset[31:0]), //i
    .io_fetchGroupIn_payload_predecodeInfos_3_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isIdle          ), //i
    .io_fetchGroupIn_payload_branchMask                    (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_branchMask[3:0]                  ), //i
    .io_fetchGroupIn_payload_fault                         (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_fault                            ), //i
    .io_fetchGroupIn_payload_numValidInstructions          (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_numValidInstructions[2:0]        ), //i
    .io_fetchGroupIn_payload_startInstructionIndex         (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_startInstructionIndex[1:0]       ), //i
    .io_bpuRsp_valid                                       (BpuPipelinePlugin_responseFlowOut_valid                                                             ), //i
    .io_bpuRsp_payload_isTaken                             (BpuPipelinePlugin_responseFlowOut_payload_isTaken                                                   ), //i
    .io_bpuRsp_payload_target                              (BpuPipelinePlugin_responseFlowOut_payload_target[31:0]                                              ), //i
    .io_bpuRsp_payload_transactionId                       (BpuPipelinePlugin_responseFlowOut_payload_transactionId[2:0]                                        ), //i
    .io_bpuRsp_payload_qPc                                 (BpuPipelinePlugin_responseFlowOut_payload_qPc[31:0]                                                 ), //i
    .io_fetchOutput_valid                                  (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_valid                                           ), //o
    .io_fetchOutput_ready                                  (FetchPipelinePlugin_setup_fetchOutput_io_push_ready                                                 ), //i
    .io_fetchOutput_payload_pc                             (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_pc[31:0]                                ), //o
    .io_fetchOutput_payload_instruction                    (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_instruction[31:0]                       ), //o
    .io_fetchOutput_payload_predecode_isBranch             (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isBranch                      ), //o
    .io_fetchOutput_payload_predecode_isJump               (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isJump                        ), //o
    .io_fetchOutput_payload_predecode_isDirectJump         (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isDirectJump                  ), //o
    .io_fetchOutput_payload_predecode_jumpOffset           (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_jumpOffset[31:0]              ), //o
    .io_fetchOutput_payload_predecode_isIdle               (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_predecode_isIdle                        ), //o
    .io_fetchOutput_payload_bpuPrediction_isTaken          (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_isTaken                   ), //o
    .io_fetchOutput_payload_bpuPrediction_target           (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_target[31:0]              ), //o
    .io_fetchOutput_payload_bpuPrediction_wasPredicted     (FetchPipelinePlugin_logic_dispatcher_io_fetchOutput_payload_bpuPrediction_wasPredicted              ), //o
    .io_bpuQuery_valid                                     (FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_valid                                              ), //o
    .io_bpuQuery_payload_pc                                (FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_payload_pc[31:0]                                   ), //o
    .io_bpuQuery_payload_transactionId                     (FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_payload_transactionId[2:0]                         ), //o
    .io_softRedirect_valid                                 (FetchPipelinePlugin_logic_dispatcher_io_softRedirect_valid                                          ), //o
    .io_softRedirect_payload                               (FetchPipelinePlugin_logic_dispatcher_io_softRedirect_payload[31:0]                                  ), //o
    .io_flush                                              (FetchPipelinePlugin_logic_hardRedirect_valid                                                        ), //i
    .clk                                                   (clk                                                                                                 ), //i
    .reset                                                 (reset                                                                                               )  //i
  );
  StreamFifo_12 FetchPipelinePlugin_logic_s4_logic_predecodedGroups (
    .io_push_valid                                 (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_valid                                    ), //i
    .io_push_ready                                 (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_ready                                    ), //o
    .io_push_payload_pc                            (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_pc[31:0]                         ), //i
    .io_push_payload_instructions_0                (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_0[31:0]             ), //i
    .io_push_payload_instructions_1                (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_1[31:0]             ), //i
    .io_push_payload_instructions_2                (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_2[31:0]             ), //i
    .io_push_payload_instructions_3                (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_3[31:0]             ), //i
    .io_push_payload_predecodeInfos_0_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isBranch        ), //i
    .io_push_payload_predecodeInfos_0_isJump       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isJump          ), //i
    .io_push_payload_predecodeInfos_0_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isDirectJump    ), //i
    .io_push_payload_predecodeInfos_0_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_jumpOffset[31:0]), //i
    .io_push_payload_predecodeInfos_0_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isIdle          ), //i
    .io_push_payload_predecodeInfos_1_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isBranch        ), //i
    .io_push_payload_predecodeInfos_1_isJump       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isJump          ), //i
    .io_push_payload_predecodeInfos_1_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isDirectJump    ), //i
    .io_push_payload_predecodeInfos_1_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_jumpOffset[31:0]), //i
    .io_push_payload_predecodeInfos_1_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isIdle          ), //i
    .io_push_payload_predecodeInfos_2_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isBranch        ), //i
    .io_push_payload_predecodeInfos_2_isJump       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isJump          ), //i
    .io_push_payload_predecodeInfos_2_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isDirectJump    ), //i
    .io_push_payload_predecodeInfos_2_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_jumpOffset[31:0]), //i
    .io_push_payload_predecodeInfos_2_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isIdle          ), //i
    .io_push_payload_predecodeInfos_3_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isBranch        ), //i
    .io_push_payload_predecodeInfos_3_isJump       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isJump          ), //i
    .io_push_payload_predecodeInfos_3_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isDirectJump    ), //i
    .io_push_payload_predecodeInfos_3_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_jumpOffset[31:0]), //i
    .io_push_payload_predecodeInfos_3_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isIdle          ), //i
    .io_push_payload_branchMask                    (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_branchMask[3:0]                  ), //i
    .io_push_payload_fault                         (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_fault                            ), //i
    .io_push_payload_numValidInstructions          (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_numValidInstructions[2:0]        ), //i
    .io_push_payload_startInstructionIndex         (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_startInstructionIndex[1:0]       ), //i
    .io_pop_valid                                  (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_valid                                     ), //o
    .io_pop_ready                                  (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_ready                                     ), //i
    .io_pop_payload_pc                             (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_pc[31:0]                          ), //o
    .io_pop_payload_instructions_0                 (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_0[31:0]              ), //o
    .io_pop_payload_instructions_1                 (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_1[31:0]              ), //o
    .io_pop_payload_instructions_2                 (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_2[31:0]              ), //o
    .io_pop_payload_instructions_3                 (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_instructions_3[31:0]              ), //o
    .io_pop_payload_predecodeInfos_0_isBranch      (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isBranch         ), //o
    .io_pop_payload_predecodeInfos_0_isJump        (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isJump           ), //o
    .io_pop_payload_predecodeInfos_0_isDirectJump  (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isDirectJump     ), //o
    .io_pop_payload_predecodeInfos_0_jumpOffset    (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_jumpOffset[31:0] ), //o
    .io_pop_payload_predecodeInfos_0_isIdle        (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isIdle           ), //o
    .io_pop_payload_predecodeInfos_1_isBranch      (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isBranch         ), //o
    .io_pop_payload_predecodeInfos_1_isJump        (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isJump           ), //o
    .io_pop_payload_predecodeInfos_1_isDirectJump  (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isDirectJump     ), //o
    .io_pop_payload_predecodeInfos_1_jumpOffset    (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_jumpOffset[31:0] ), //o
    .io_pop_payload_predecodeInfos_1_isIdle        (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isIdle           ), //o
    .io_pop_payload_predecodeInfos_2_isBranch      (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isBranch         ), //o
    .io_pop_payload_predecodeInfos_2_isJump        (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isJump           ), //o
    .io_pop_payload_predecodeInfos_2_isDirectJump  (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isDirectJump     ), //o
    .io_pop_payload_predecodeInfos_2_jumpOffset    (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_jumpOffset[31:0] ), //o
    .io_pop_payload_predecodeInfos_2_isIdle        (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isIdle           ), //o
    .io_pop_payload_predecodeInfos_3_isBranch      (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isBranch         ), //o
    .io_pop_payload_predecodeInfos_3_isJump        (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isJump           ), //o
    .io_pop_payload_predecodeInfos_3_isDirectJump  (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isDirectJump     ), //o
    .io_pop_payload_predecodeInfos_3_jumpOffset    (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_jumpOffset[31:0] ), //o
    .io_pop_payload_predecodeInfos_3_isIdle        (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isIdle           ), //o
    .io_pop_payload_branchMask                     (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_branchMask[3:0]                   ), //o
    .io_pop_payload_fault                          (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_fault                             ), //o
    .io_pop_payload_numValidInstructions           (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_numValidInstructions[2:0]         ), //o
    .io_pop_payload_startInstructionIndex          (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_startInstructionIndex[1:0]        ), //o
    .io_flush                                      (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_flush                                         ), //i
    .io_occupancy                                  (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_occupancy[1:0]                                ), //o
    .io_availability                               (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_availability[1:0]                             ), //o
    .clk                                           (clk                                                                                                  ), //i
    .reset                                         (reset                                                                                                )  //i
  );
  InstructionPredecoder FetchPipelinePlugin_logic_s4_logic_predecoders_0 (
    .io_instruction                (FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_instruction[31:0]             ), //i
    .io_predecodeInfo_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isBranch        ), //o
    .io_predecodeInfo_isJump       (FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isJump          ), //o
    .io_predecodeInfo_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isDirectJump    ), //o
    .io_predecodeInfo_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_jumpOffset[31:0]), //o
    .io_predecodeInfo_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isIdle          ), //o
    .clk                           (clk                                                                               ), //i
    .reset                         (reset                                                                             )  //i
  );
  InstructionPredecoder FetchPipelinePlugin_logic_s4_logic_predecoders_1 (
    .io_instruction                (FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_instruction[31:0]             ), //i
    .io_predecodeInfo_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isBranch        ), //o
    .io_predecodeInfo_isJump       (FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isJump          ), //o
    .io_predecodeInfo_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isDirectJump    ), //o
    .io_predecodeInfo_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_jumpOffset[31:0]), //o
    .io_predecodeInfo_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isIdle          ), //o
    .clk                           (clk                                                                               ), //i
    .reset                         (reset                                                                             )  //i
  );
  InstructionPredecoder FetchPipelinePlugin_logic_s4_logic_predecoders_2 (
    .io_instruction                (FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_instruction[31:0]             ), //i
    .io_predecodeInfo_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isBranch        ), //o
    .io_predecodeInfo_isJump       (FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isJump          ), //o
    .io_predecodeInfo_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isDirectJump    ), //o
    .io_predecodeInfo_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_jumpOffset[31:0]), //o
    .io_predecodeInfo_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isIdle          ), //o
    .clk                           (clk                                                                               ), //i
    .reset                         (reset                                                                             )  //i
  );
  InstructionPredecoder FetchPipelinePlugin_logic_s4_logic_predecoders_3 (
    .io_instruction                (FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_instruction[31:0]             ), //i
    .io_predecodeInfo_isBranch     (FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isBranch        ), //o
    .io_predecodeInfo_isJump       (FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isJump          ), //o
    .io_predecodeInfo_isDirectJump (FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isDirectJump    ), //o
    .io_predecodeInfo_jumpOffset   (FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_jumpOffset[31:0]), //o
    .io_predecodeInfo_isIdle       (FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isIdle          ), //o
    .clk                           (clk                                                                               ), //i
    .reset                         (reset                                                                             )  //i
  );
  SplitGmbToAxi4Bridge CoreMemSysPlugin_logic_readBridges_0 (
    .io_gmbIn_read_cmd_valid                (_zz_LoadQueuePlugin_logic_loadQueue_mmioCmdFired                         ), //i
    .io_gmbIn_read_cmd_ready                (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_cmd_ready             ), //o
    .io_gmbIn_read_cmd_payload_address      (LoadQueuePlugin_logic_loadQueue_slots_0_address[31:0]                    ), //i
    .io_gmbIn_read_cmd_payload_id           (LoadQueuePlugin_logic_loadQueue_slots_0_robPtr[3:0]                      ), //i
    .io_gmbIn_read_rsp_valid                (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_valid             ), //o
    .io_gmbIn_read_rsp_ready                (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_ready             ), //i
    .io_gmbIn_read_rsp_payload_data         (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_payload_data[31:0]), //o
    .io_gmbIn_read_rsp_payload_error        (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_payload_error     ), //o
    .io_gmbIn_read_rsp_payload_id           (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_payload_id[3:0]   ), //o
    .io_gmbIn_write_cmd_valid               (1'b0                                                                     ), //i
    .io_gmbIn_write_cmd_ready               (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_write_cmd_ready            ), //o
    .io_gmbIn_write_cmd_payload_address     (32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx                                     ), //i
    .io_gmbIn_write_cmd_payload_data        (32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx                                     ), //i
    .io_gmbIn_write_cmd_payload_byteEnables (4'bxxxx                                                                  ), //i
    .io_gmbIn_write_cmd_payload_id          (4'bxxxx                                                                  ), //i
    .io_gmbIn_write_cmd_payload_last        (1'bx                                                                     ), //i
    .io_gmbIn_write_rsp_valid               (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_write_rsp_valid            ), //o
    .io_gmbIn_write_rsp_ready               (1'b1                                                                     ), //i
    .io_gmbIn_write_rsp_payload_error       (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_write_rsp_payload_error    ), //o
    .io_gmbIn_write_rsp_payload_id          (CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_write_rsp_payload_id[3:0]  ), //o
    .io_axiOut_aw_valid                     (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_valid                  ), //o
    .io_axiOut_aw_ready                     (io_axiOut_writeOnly_aw_ready_1                                           ), //i
    .io_axiOut_aw_payload_addr              (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_addr[31:0]     ), //o
    .io_axiOut_aw_payload_id                (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_id[3:0]        ), //o
    .io_axiOut_aw_payload_len               (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_len[7:0]       ), //o
    .io_axiOut_aw_payload_size              (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_size[2:0]      ), //o
    .io_axiOut_aw_payload_burst             (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_burst[1:0]     ), //o
    .io_axiOut_w_valid                      (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_valid                   ), //o
    .io_axiOut_w_ready                      (io_axiOut_writeOnly_w_ready_1                                            ), //i
    .io_axiOut_w_payload_data               (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_data[31:0]      ), //o
    .io_axiOut_w_payload_strb               (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_strb[3:0]       ), //o
    .io_axiOut_w_payload_last               (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_last            ), //o
    .io_axiOut_b_valid                      (io_axiOut_writeOnly_b_valid_1                                            ), //i
    .io_axiOut_b_ready                      (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_b_ready                   ), //o
    .io_axiOut_b_payload_id                 (io_axiOut_writeOnly_b_payload_id_1[3:0]                                  ), //i
    .io_axiOut_b_payload_resp               (io_axiOut_writeOnly_b_payload_resp_1[1:0]                                ), //i
    .io_axiOut_ar_valid                     (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_valid                  ), //o
    .io_axiOut_ar_ready                     (io_axiOut_readOnly_ar_ready_1                                            ), //i
    .io_axiOut_ar_payload_addr              (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_addr[31:0]     ), //o
    .io_axiOut_ar_payload_id                (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_id[3:0]        ), //o
    .io_axiOut_ar_payload_len               (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_len[7:0]       ), //o
    .io_axiOut_ar_payload_size              (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_size[2:0]      ), //o
    .io_axiOut_ar_payload_burst             (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_burst[1:0]     ), //o
    .io_axiOut_r_valid                      (io_axiOut_readOnly_r_valid_1                                             ), //i
    .io_axiOut_r_ready                      (CoreMemSysPlugin_logic_readBridges_0_io_axiOut_r_ready                   ), //o
    .io_axiOut_r_payload_data               (io_axiOut_readOnly_r_payload_data_1[31:0]                                ), //i
    .io_axiOut_r_payload_id                 (io_axiOut_readOnly_r_payload_id_1[3:0]                                   ), //i
    .io_axiOut_r_payload_resp               (io_axiOut_readOnly_r_payload_resp_1[1:0]                                 ), //i
    .io_axiOut_r_payload_last               (io_axiOut_readOnly_r_payload_last_1                                      ), //i
    .clk                                    (clk                                                                      ), //i
    .reset                                  (reset                                                                    )  //i
  );
  SplitGmbToAxi4Bridge CoreMemSysPlugin_logic_writeBridges_0 (
    .io_gmbIn_read_cmd_valid                (1'b0                                                                      ), //i
    .io_gmbIn_read_cmd_ready                (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_cmd_ready             ), //o
    .io_gmbIn_read_cmd_payload_address      (32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx                                      ), //i
    .io_gmbIn_read_cmd_payload_id           (4'bxxxx                                                                   ), //i
    .io_gmbIn_read_rsp_valid                (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_rsp_valid             ), //o
    .io_gmbIn_read_rsp_ready                (1'b1                                                                      ), //i
    .io_gmbIn_read_rsp_payload_data         (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_rsp_payload_data[31:0]), //o
    .io_gmbIn_read_rsp_payload_error        (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_rsp_payload_error     ), //o
    .io_gmbIn_read_rsp_payload_id           (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_read_rsp_payload_id[3:0]   ), //o
    .io_gmbIn_write_cmd_valid               (StoreBufferPlugin_logic_canPopMMIOOp                                      ), //i
    .io_gmbIn_write_cmd_ready               (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_cmd_ready            ), //o
    .io_gmbIn_write_cmd_payload_address     (StoreBufferPlugin_logic_slots_0_addr[31:0]                                ), //i
    .io_gmbIn_write_cmd_payload_data        (StoreBufferPlugin_logic_slots_0_data[31:0]                                ), //i
    .io_gmbIn_write_cmd_payload_byteEnables (StoreBufferPlugin_logic_slots_0_be[3:0]                                   ), //i
    .io_gmbIn_write_cmd_payload_id          (StoreBufferPlugin_logic_slots_0_robPtr[3:0]                               ), //i
    .io_gmbIn_write_cmd_payload_last        (1'b1                                                                      ), //i
    .io_gmbIn_write_rsp_valid               (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_valid            ), //o
    .io_gmbIn_write_rsp_ready               (StoreBufferPlugin_logic_mmioResponseForHead                               ), //i
    .io_gmbIn_write_rsp_payload_error       (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_payload_error    ), //o
    .io_gmbIn_write_rsp_payload_id          (CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_payload_id[3:0]  ), //o
    .io_axiOut_aw_valid                     (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_valid                  ), //o
    .io_axiOut_aw_ready                     (io_axiOut_writeOnly_aw_ready                                              ), //i
    .io_axiOut_aw_payload_addr              (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_addr[31:0]     ), //o
    .io_axiOut_aw_payload_id                (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_id[3:0]        ), //o
    .io_axiOut_aw_payload_len               (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_len[7:0]       ), //o
    .io_axiOut_aw_payload_size              (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_size[2:0]      ), //o
    .io_axiOut_aw_payload_burst             (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_burst[1:0]     ), //o
    .io_axiOut_w_valid                      (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_valid                   ), //o
    .io_axiOut_w_ready                      (io_axiOut_writeOnly_w_ready                                               ), //i
    .io_axiOut_w_payload_data               (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_data[31:0]      ), //o
    .io_axiOut_w_payload_strb               (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_strb[3:0]       ), //o
    .io_axiOut_w_payload_last               (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_last            ), //o
    .io_axiOut_b_valid                      (io_axiOut_writeOnly_b_valid                                               ), //i
    .io_axiOut_b_ready                      (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_b_ready                   ), //o
    .io_axiOut_b_payload_id                 (io_axiOut_writeOnly_b_payload_id[3:0]                                     ), //i
    .io_axiOut_b_payload_resp               (io_axiOut_writeOnly_b_payload_resp[1:0]                                   ), //i
    .io_axiOut_ar_valid                     (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_valid                  ), //o
    .io_axiOut_ar_ready                     (io_axiOut_readOnly_ar_ready                                               ), //i
    .io_axiOut_ar_payload_addr              (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_addr[31:0]     ), //o
    .io_axiOut_ar_payload_id                (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_id[3:0]        ), //o
    .io_axiOut_ar_payload_len               (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_len[7:0]       ), //o
    .io_axiOut_ar_payload_size              (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_size[2:0]      ), //o
    .io_axiOut_ar_payload_burst             (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_burst[1:0]     ), //o
    .io_axiOut_r_valid                      (io_axiOut_readOnly_r_valid                                                ), //i
    .io_axiOut_r_ready                      (CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_r_ready                   ), //o
    .io_axiOut_r_payload_data               (io_axiOut_readOnly_r_payload_data[31:0]                                   ), //i
    .io_axiOut_r_payload_id                 (io_axiOut_readOnly_r_payload_id[3:0]                                      ), //i
    .io_axiOut_r_payload_resp               (io_axiOut_readOnly_r_payload_resp[1:0]                                    ), //i
    .io_axiOut_r_payload_last               (io_axiOut_readOnly_r_payload_last                                         ), //i
    .clk                                    (clk                                                                       ), //i
    .reset                                  (reset                                                                     )  //i
  );
  Axi4ReadOnlyDecoder io_axiOut_readOnly_decoder (
    .io_input_ar_valid             (io_axiOut_readOnly_ar_valid                                  ), //i
    .io_input_ar_ready             (io_axiOut_readOnly_decoder_io_input_ar_ready                 ), //o
    .io_input_ar_payload_addr      (io_axiOut_readOnly_ar_payload_addr[31:0]                     ), //i
    .io_input_ar_payload_id        (io_axiOut_readOnly_ar_payload_id[3:0]                        ), //i
    .io_input_ar_payload_len       (io_axiOut_readOnly_ar_payload_len[7:0]                       ), //i
    .io_input_ar_payload_size      (io_axiOut_readOnly_ar_payload_size[2:0]                      ), //i
    .io_input_ar_payload_burst     (io_axiOut_readOnly_ar_payload_burst[1:0]                     ), //i
    .io_input_r_valid              (io_axiOut_readOnly_decoder_io_input_r_valid                  ), //o
    .io_input_r_ready              (io_axiOut_readOnly_r_ready                                   ), //i
    .io_input_r_payload_data       (io_axiOut_readOnly_decoder_io_input_r_payload_data[31:0]     ), //o
    .io_input_r_payload_id         (io_axiOut_readOnly_decoder_io_input_r_payload_id[3:0]        ), //o
    .io_input_r_payload_resp       (io_axiOut_readOnly_decoder_io_input_r_payload_resp[1:0]      ), //o
    .io_input_r_payload_last       (io_axiOut_readOnly_decoder_io_input_r_payload_last           ), //o
    .io_outputs_0_ar_valid         (io_axiOut_readOnly_decoder_io_outputs_0_ar_valid             ), //o
    .io_outputs_0_ar_ready         (io_outputs_0_ar_validPipe_fire                               ), //i
    .io_outputs_0_ar_payload_addr  (io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_addr[31:0]), //o
    .io_outputs_0_ar_payload_id    (io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_id[3:0]   ), //o
    .io_outputs_0_ar_payload_len   (io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_len[7:0]  ), //o
    .io_outputs_0_ar_payload_size  (io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_size[2:0] ), //o
    .io_outputs_0_ar_payload_burst (io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_burst[1:0]), //o
    .io_outputs_0_r_valid          (axi4ReadOnlyArbiter_3_io_inputs_0_r_valid                    ), //i
    .io_outputs_0_r_ready          (io_axiOut_readOnly_decoder_io_outputs_0_r_ready              ), //o
    .io_outputs_0_r_payload_data   (axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_data[31:0]       ), //i
    .io_outputs_0_r_payload_id     (io_axiOut_readOnly_decoder_io_outputs_0_r_payload_id[3:0]    ), //i
    .io_outputs_0_r_payload_resp   (axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_resp[1:0]        ), //i
    .io_outputs_0_r_payload_last   (axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_last             ), //i
    .io_outputs_1_ar_valid         (io_axiOut_readOnly_decoder_io_outputs_1_ar_valid             ), //o
    .io_outputs_1_ar_ready         (io_outputs_1_ar_validPipe_fire                               ), //i
    .io_outputs_1_ar_payload_addr  (io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_addr[31:0]), //o
    .io_outputs_1_ar_payload_id    (io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_id[3:0]   ), //o
    .io_outputs_1_ar_payload_len   (io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_len[7:0]  ), //o
    .io_outputs_1_ar_payload_size  (io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_size[2:0] ), //o
    .io_outputs_1_ar_payload_burst (io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_burst[1:0]), //o
    .io_outputs_1_r_valid          (axi4ReadOnlyArbiter_4_io_inputs_0_r_valid                    ), //i
    .io_outputs_1_r_ready          (io_axiOut_readOnly_decoder_io_outputs_1_r_ready              ), //o
    .io_outputs_1_r_payload_data   (axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_data[31:0]       ), //i
    .io_outputs_1_r_payload_id     (io_axiOut_readOnly_decoder_io_outputs_1_r_payload_id[3:0]    ), //i
    .io_outputs_1_r_payload_resp   (axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_resp[1:0]        ), //i
    .io_outputs_1_r_payload_last   (axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_last             ), //i
    .io_outputs_2_ar_valid         (io_axiOut_readOnly_decoder_io_outputs_2_ar_valid             ), //o
    .io_outputs_2_ar_ready         (io_outputs_2_ar_validPipe_fire                               ), //i
    .io_outputs_2_ar_payload_addr  (io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_addr[31:0]), //o
    .io_outputs_2_ar_payload_id    (io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_id[3:0]   ), //o
    .io_outputs_2_ar_payload_len   (io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_len[7:0]  ), //o
    .io_outputs_2_ar_payload_size  (io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_size[2:0] ), //o
    .io_outputs_2_ar_payload_burst (io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_burst[1:0]), //o
    .io_outputs_2_r_valid          (axi4ReadOnlyArbiter_5_io_inputs_0_r_valid                    ), //i
    .io_outputs_2_r_ready          (io_axiOut_readOnly_decoder_io_outputs_2_r_ready              ), //o
    .io_outputs_2_r_payload_data   (axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_data[31:0]       ), //i
    .io_outputs_2_r_payload_id     (io_axiOut_readOnly_decoder_io_outputs_2_r_payload_id[3:0]    ), //i
    .io_outputs_2_r_payload_resp   (axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_resp[1:0]        ), //i
    .io_outputs_2_r_payload_last   (axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_last             ), //i
    .clk                           (clk                                                          ), //i
    .reset                         (reset                                                        )  //i
  );
  Axi4WriteOnlyDecoder io_axiOut_writeOnly_decoder (
    .io_input_aw_valid             (io_axiOut_writeOnly_aw_valid                                  ), //i
    .io_input_aw_ready             (io_axiOut_writeOnly_decoder_io_input_aw_ready                 ), //o
    .io_input_aw_payload_addr      (io_axiOut_writeOnly_aw_payload_addr[31:0]                     ), //i
    .io_input_aw_payload_id        (io_axiOut_writeOnly_aw_payload_id[3:0]                        ), //i
    .io_input_aw_payload_len       (io_axiOut_writeOnly_aw_payload_len[7:0]                       ), //i
    .io_input_aw_payload_size      (io_axiOut_writeOnly_aw_payload_size[2:0]                      ), //i
    .io_input_aw_payload_burst     (io_axiOut_writeOnly_aw_payload_burst[1:0]                     ), //i
    .io_input_w_valid              (io_axiOut_writeOnly_w_valid                                   ), //i
    .io_input_w_ready              (io_axiOut_writeOnly_decoder_io_input_w_ready                  ), //o
    .io_input_w_payload_data       (io_axiOut_writeOnly_w_payload_data[31:0]                      ), //i
    .io_input_w_payload_strb       (io_axiOut_writeOnly_w_payload_strb[3:0]                       ), //i
    .io_input_w_payload_last       (io_axiOut_writeOnly_w_payload_last                            ), //i
    .io_input_b_valid              (io_axiOut_writeOnly_decoder_io_input_b_valid                  ), //o
    .io_input_b_ready              (io_axiOut_writeOnly_b_ready                                   ), //i
    .io_input_b_payload_id         (io_axiOut_writeOnly_decoder_io_input_b_payload_id[3:0]        ), //o
    .io_input_b_payload_resp       (io_axiOut_writeOnly_decoder_io_input_b_payload_resp[1:0]      ), //o
    .io_outputs_0_aw_valid         (io_axiOut_writeOnly_decoder_io_outputs_0_aw_valid             ), //o
    .io_outputs_0_aw_ready         (io_outputs_0_aw_validPipe_fire                                ), //i
    .io_outputs_0_aw_payload_addr  (io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_addr[31:0]), //o
    .io_outputs_0_aw_payload_id    (io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_id[3:0]   ), //o
    .io_outputs_0_aw_payload_len   (io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_len[7:0]  ), //o
    .io_outputs_0_aw_payload_size  (io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_size[2:0] ), //o
    .io_outputs_0_aw_payload_burst (io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_burst[1:0]), //o
    .io_outputs_0_w_valid          (io_axiOut_writeOnly_decoder_io_outputs_0_w_valid              ), //o
    .io_outputs_0_w_ready          (axi4WriteOnlyArbiter_3_io_inputs_0_w_ready                    ), //i
    .io_outputs_0_w_payload_data   (io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_data[31:0] ), //o
    .io_outputs_0_w_payload_strb   (io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]  ), //o
    .io_outputs_0_w_payload_last   (io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_last       ), //o
    .io_outputs_0_b_valid          (axi4WriteOnlyArbiter_3_io_inputs_0_b_valid                    ), //i
    .io_outputs_0_b_ready          (io_axiOut_writeOnly_decoder_io_outputs_0_b_ready              ), //o
    .io_outputs_0_b_payload_id     (io_axiOut_writeOnly_decoder_io_outputs_0_b_payload_id[3:0]    ), //i
    .io_outputs_0_b_payload_resp   (axi4WriteOnlyArbiter_3_io_inputs_0_b_payload_resp[1:0]        ), //i
    .io_outputs_1_aw_valid         (io_axiOut_writeOnly_decoder_io_outputs_1_aw_valid             ), //o
    .io_outputs_1_aw_ready         (io_outputs_1_aw_validPipe_fire                                ), //i
    .io_outputs_1_aw_payload_addr  (io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_addr[31:0]), //o
    .io_outputs_1_aw_payload_id    (io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_id[3:0]   ), //o
    .io_outputs_1_aw_payload_len   (io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_len[7:0]  ), //o
    .io_outputs_1_aw_payload_size  (io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_size[2:0] ), //o
    .io_outputs_1_aw_payload_burst (io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_burst[1:0]), //o
    .io_outputs_1_w_valid          (io_axiOut_writeOnly_decoder_io_outputs_1_w_valid              ), //o
    .io_outputs_1_w_ready          (axi4WriteOnlyArbiter_4_io_inputs_0_w_ready                    ), //i
    .io_outputs_1_w_payload_data   (io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_data[31:0] ), //o
    .io_outputs_1_w_payload_strb   (io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_strb[3:0]  ), //o
    .io_outputs_1_w_payload_last   (io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_last       ), //o
    .io_outputs_1_b_valid          (axi4WriteOnlyArbiter_4_io_inputs_0_b_valid                    ), //i
    .io_outputs_1_b_ready          (io_axiOut_writeOnly_decoder_io_outputs_1_b_ready              ), //o
    .io_outputs_1_b_payload_id     (io_axiOut_writeOnly_decoder_io_outputs_1_b_payload_id[3:0]    ), //i
    .io_outputs_1_b_payload_resp   (axi4WriteOnlyArbiter_4_io_inputs_0_b_payload_resp[1:0]        ), //i
    .io_outputs_2_aw_valid         (io_axiOut_writeOnly_decoder_io_outputs_2_aw_valid             ), //o
    .io_outputs_2_aw_ready         (io_outputs_2_aw_validPipe_fire                                ), //i
    .io_outputs_2_aw_payload_addr  (io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_addr[31:0]), //o
    .io_outputs_2_aw_payload_id    (io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_id[3:0]   ), //o
    .io_outputs_2_aw_payload_len   (io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_len[7:0]  ), //o
    .io_outputs_2_aw_payload_size  (io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_size[2:0] ), //o
    .io_outputs_2_aw_payload_burst (io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_burst[1:0]), //o
    .io_outputs_2_w_valid          (io_axiOut_writeOnly_decoder_io_outputs_2_w_valid              ), //o
    .io_outputs_2_w_ready          (axi4WriteOnlyArbiter_5_io_inputs_0_w_ready                    ), //i
    .io_outputs_2_w_payload_data   (io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_data[31:0] ), //o
    .io_outputs_2_w_payload_strb   (io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_strb[3:0]  ), //o
    .io_outputs_2_w_payload_last   (io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_last       ), //o
    .io_outputs_2_b_valid          (axi4WriteOnlyArbiter_5_io_inputs_0_b_valid                    ), //i
    .io_outputs_2_b_ready          (io_axiOut_writeOnly_decoder_io_outputs_2_b_ready              ), //o
    .io_outputs_2_b_payload_id     (io_axiOut_writeOnly_decoder_io_outputs_2_b_payload_id[3:0]    ), //i
    .io_outputs_2_b_payload_resp   (axi4WriteOnlyArbiter_5_io_inputs_0_b_payload_resp[1:0]        ), //i
    .clk                           (clk                                                           ), //i
    .reset                         (reset                                                         )  //i
  );
  Axi4ReadOnlyDecoder io_axiOut_readOnly_decoder_1 (
    .io_input_ar_valid             (io_axiOut_readOnly_ar_valid_1                                  ), //i
    .io_input_ar_ready             (io_axiOut_readOnly_decoder_1_io_input_ar_ready                 ), //o
    .io_input_ar_payload_addr      (io_axiOut_readOnly_ar_payload_addr_1[31:0]                     ), //i
    .io_input_ar_payload_id        (io_axiOut_readOnly_ar_payload_id_1[3:0]                        ), //i
    .io_input_ar_payload_len       (io_axiOut_readOnly_ar_payload_len_1[7:0]                       ), //i
    .io_input_ar_payload_size      (io_axiOut_readOnly_ar_payload_size_1[2:0]                      ), //i
    .io_input_ar_payload_burst     (io_axiOut_readOnly_ar_payload_burst_1[1:0]                     ), //i
    .io_input_r_valid              (io_axiOut_readOnly_decoder_1_io_input_r_valid                  ), //o
    .io_input_r_ready              (io_axiOut_readOnly_r_ready_1                                   ), //i
    .io_input_r_payload_data       (io_axiOut_readOnly_decoder_1_io_input_r_payload_data[31:0]     ), //o
    .io_input_r_payload_id         (io_axiOut_readOnly_decoder_1_io_input_r_payload_id[3:0]        ), //o
    .io_input_r_payload_resp       (io_axiOut_readOnly_decoder_1_io_input_r_payload_resp[1:0]      ), //o
    .io_input_r_payload_last       (io_axiOut_readOnly_decoder_1_io_input_r_payload_last           ), //o
    .io_outputs_0_ar_valid         (io_axiOut_readOnly_decoder_1_io_outputs_0_ar_valid             ), //o
    .io_outputs_0_ar_ready         (io_outputs_0_ar_validPipe_fire_1                               ), //i
    .io_outputs_0_ar_payload_addr  (io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_addr[31:0]), //o
    .io_outputs_0_ar_payload_id    (io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_id[3:0]   ), //o
    .io_outputs_0_ar_payload_len   (io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_len[7:0]  ), //o
    .io_outputs_0_ar_payload_size  (io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_size[2:0] ), //o
    .io_outputs_0_ar_payload_burst (io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_burst[1:0]), //o
    .io_outputs_0_r_valid          (axi4ReadOnlyArbiter_3_io_inputs_1_r_valid                      ), //i
    .io_outputs_0_r_ready          (io_axiOut_readOnly_decoder_1_io_outputs_0_r_ready              ), //o
    .io_outputs_0_r_payload_data   (axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_data[31:0]         ), //i
    .io_outputs_0_r_payload_id     (io_axiOut_readOnly_decoder_1_io_outputs_0_r_payload_id[3:0]    ), //i
    .io_outputs_0_r_payload_resp   (axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_resp[1:0]          ), //i
    .io_outputs_0_r_payload_last   (axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_last               ), //i
    .io_outputs_1_ar_valid         (io_axiOut_readOnly_decoder_1_io_outputs_1_ar_valid             ), //o
    .io_outputs_1_ar_ready         (io_outputs_1_ar_validPipe_fire_1                               ), //i
    .io_outputs_1_ar_payload_addr  (io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_addr[31:0]), //o
    .io_outputs_1_ar_payload_id    (io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_id[3:0]   ), //o
    .io_outputs_1_ar_payload_len   (io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_len[7:0]  ), //o
    .io_outputs_1_ar_payload_size  (io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_size[2:0] ), //o
    .io_outputs_1_ar_payload_burst (io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_burst[1:0]), //o
    .io_outputs_1_r_valid          (axi4ReadOnlyArbiter_4_io_inputs_1_r_valid                      ), //i
    .io_outputs_1_r_ready          (io_axiOut_readOnly_decoder_1_io_outputs_1_r_ready              ), //o
    .io_outputs_1_r_payload_data   (axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_data[31:0]         ), //i
    .io_outputs_1_r_payload_id     (io_axiOut_readOnly_decoder_1_io_outputs_1_r_payload_id[3:0]    ), //i
    .io_outputs_1_r_payload_resp   (axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_resp[1:0]          ), //i
    .io_outputs_1_r_payload_last   (axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_last               ), //i
    .io_outputs_2_ar_valid         (io_axiOut_readOnly_decoder_1_io_outputs_2_ar_valid             ), //o
    .io_outputs_2_ar_ready         (io_outputs_2_ar_validPipe_fire_1                               ), //i
    .io_outputs_2_ar_payload_addr  (io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_addr[31:0]), //o
    .io_outputs_2_ar_payload_id    (io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_id[3:0]   ), //o
    .io_outputs_2_ar_payload_len   (io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_len[7:0]  ), //o
    .io_outputs_2_ar_payload_size  (io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_size[2:0] ), //o
    .io_outputs_2_ar_payload_burst (io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_burst[1:0]), //o
    .io_outputs_2_r_valid          (axi4ReadOnlyArbiter_5_io_inputs_1_r_valid                      ), //i
    .io_outputs_2_r_ready          (io_axiOut_readOnly_decoder_1_io_outputs_2_r_ready              ), //o
    .io_outputs_2_r_payload_data   (axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_data[31:0]         ), //i
    .io_outputs_2_r_payload_id     (io_axiOut_readOnly_decoder_1_io_outputs_2_r_payload_id[3:0]    ), //i
    .io_outputs_2_r_payload_resp   (axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_resp[1:0]          ), //i
    .io_outputs_2_r_payload_last   (axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_last               ), //i
    .clk                           (clk                                                            ), //i
    .reset                         (reset                                                          )  //i
  );
  Axi4WriteOnlyDecoder io_axiOut_writeOnly_decoder_1 (
    .io_input_aw_valid             (io_axiOut_writeOnly_aw_valid_1                                  ), //i
    .io_input_aw_ready             (io_axiOut_writeOnly_decoder_1_io_input_aw_ready                 ), //o
    .io_input_aw_payload_addr      (io_axiOut_writeOnly_aw_payload_addr_1[31:0]                     ), //i
    .io_input_aw_payload_id        (io_axiOut_writeOnly_aw_payload_id_1[3:0]                        ), //i
    .io_input_aw_payload_len       (io_axiOut_writeOnly_aw_payload_len_1[7:0]                       ), //i
    .io_input_aw_payload_size      (io_axiOut_writeOnly_aw_payload_size_1[2:0]                      ), //i
    .io_input_aw_payload_burst     (io_axiOut_writeOnly_aw_payload_burst_1[1:0]                     ), //i
    .io_input_w_valid              (io_axiOut_writeOnly_w_valid_1                                   ), //i
    .io_input_w_ready              (io_axiOut_writeOnly_decoder_1_io_input_w_ready                  ), //o
    .io_input_w_payload_data       (io_axiOut_writeOnly_w_payload_data_1[31:0]                      ), //i
    .io_input_w_payload_strb       (io_axiOut_writeOnly_w_payload_strb_1[3:0]                       ), //i
    .io_input_w_payload_last       (io_axiOut_writeOnly_w_payload_last_1                            ), //i
    .io_input_b_valid              (io_axiOut_writeOnly_decoder_1_io_input_b_valid                  ), //o
    .io_input_b_ready              (io_axiOut_writeOnly_b_ready_1                                   ), //i
    .io_input_b_payload_id         (io_axiOut_writeOnly_decoder_1_io_input_b_payload_id[3:0]        ), //o
    .io_input_b_payload_resp       (io_axiOut_writeOnly_decoder_1_io_input_b_payload_resp[1:0]      ), //o
    .io_outputs_0_aw_valid         (io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_valid             ), //o
    .io_outputs_0_aw_ready         (io_outputs_0_aw_validPipe_fire_1                                ), //i
    .io_outputs_0_aw_payload_addr  (io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_addr[31:0]), //o
    .io_outputs_0_aw_payload_id    (io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_id[3:0]   ), //o
    .io_outputs_0_aw_payload_len   (io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_len[7:0]  ), //o
    .io_outputs_0_aw_payload_size  (io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_size[2:0] ), //o
    .io_outputs_0_aw_payload_burst (io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_burst[1:0]), //o
    .io_outputs_0_w_valid          (io_axiOut_writeOnly_decoder_1_io_outputs_0_w_valid              ), //o
    .io_outputs_0_w_ready          (axi4WriteOnlyArbiter_3_io_inputs_1_w_ready                      ), //i
    .io_outputs_0_w_payload_data   (io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_data[31:0] ), //o
    .io_outputs_0_w_payload_strb   (io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_strb[3:0]  ), //o
    .io_outputs_0_w_payload_last   (io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_last       ), //o
    .io_outputs_0_b_valid          (axi4WriteOnlyArbiter_3_io_inputs_1_b_valid                      ), //i
    .io_outputs_0_b_ready          (io_axiOut_writeOnly_decoder_1_io_outputs_0_b_ready              ), //o
    .io_outputs_0_b_payload_id     (io_axiOut_writeOnly_decoder_1_io_outputs_0_b_payload_id[3:0]    ), //i
    .io_outputs_0_b_payload_resp   (axi4WriteOnlyArbiter_3_io_inputs_1_b_payload_resp[1:0]          ), //i
    .io_outputs_1_aw_valid         (io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_valid             ), //o
    .io_outputs_1_aw_ready         (io_outputs_1_aw_validPipe_fire_1                                ), //i
    .io_outputs_1_aw_payload_addr  (io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_addr[31:0]), //o
    .io_outputs_1_aw_payload_id    (io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_id[3:0]   ), //o
    .io_outputs_1_aw_payload_len   (io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_len[7:0]  ), //o
    .io_outputs_1_aw_payload_size  (io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_size[2:0] ), //o
    .io_outputs_1_aw_payload_burst (io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_burst[1:0]), //o
    .io_outputs_1_w_valid          (io_axiOut_writeOnly_decoder_1_io_outputs_1_w_valid              ), //o
    .io_outputs_1_w_ready          (axi4WriteOnlyArbiter_4_io_inputs_1_w_ready                      ), //i
    .io_outputs_1_w_payload_data   (io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_data[31:0] ), //o
    .io_outputs_1_w_payload_strb   (io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_strb[3:0]  ), //o
    .io_outputs_1_w_payload_last   (io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_last       ), //o
    .io_outputs_1_b_valid          (axi4WriteOnlyArbiter_4_io_inputs_1_b_valid                      ), //i
    .io_outputs_1_b_ready          (io_axiOut_writeOnly_decoder_1_io_outputs_1_b_ready              ), //o
    .io_outputs_1_b_payload_id     (io_axiOut_writeOnly_decoder_1_io_outputs_1_b_payload_id[3:0]    ), //i
    .io_outputs_1_b_payload_resp   (axi4WriteOnlyArbiter_4_io_inputs_1_b_payload_resp[1:0]          ), //i
    .io_outputs_2_aw_valid         (io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_valid             ), //o
    .io_outputs_2_aw_ready         (io_outputs_2_aw_validPipe_fire_1                                ), //i
    .io_outputs_2_aw_payload_addr  (io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_addr[31:0]), //o
    .io_outputs_2_aw_payload_id    (io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_id[3:0]   ), //o
    .io_outputs_2_aw_payload_len   (io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_len[7:0]  ), //o
    .io_outputs_2_aw_payload_size  (io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_size[2:0] ), //o
    .io_outputs_2_aw_payload_burst (io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_burst[1:0]), //o
    .io_outputs_2_w_valid          (io_axiOut_writeOnly_decoder_1_io_outputs_2_w_valid              ), //o
    .io_outputs_2_w_ready          (axi4WriteOnlyArbiter_5_io_inputs_1_w_ready                      ), //i
    .io_outputs_2_w_payload_data   (io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_data[31:0] ), //o
    .io_outputs_2_w_payload_strb   (io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_strb[3:0]  ), //o
    .io_outputs_2_w_payload_last   (io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_last       ), //o
    .io_outputs_2_b_valid          (axi4WriteOnlyArbiter_5_io_inputs_1_b_valid                      ), //i
    .io_outputs_2_b_ready          (io_axiOut_writeOnly_decoder_1_io_outputs_2_b_ready              ), //o
    .io_outputs_2_b_payload_id     (io_axiOut_writeOnly_decoder_1_io_outputs_2_b_payload_id[3:0]    ), //i
    .io_outputs_2_b_payload_resp   (axi4WriteOnlyArbiter_5_io_inputs_1_b_payload_resp[1:0]          ), //i
    .clk                           (clk                                                             ), //i
    .reset                         (reset                                                           )  //i
  );
  Axi4ReadOnlyDecoder_2 DataCachePlugin_setup_dcacheMaster_readOnly_decoder (
    .io_input_ar_valid             (DataCachePlugin_setup_dcacheMaster_readOnly_ar_valid                                  ), //i
    .io_input_ar_ready             (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_ar_ready                 ), //o
    .io_input_ar_payload_addr      (DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_addr[31:0]                     ), //i
    .io_input_ar_payload_id        (DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_id[2:0]                        ), //i
    .io_input_ar_payload_len       (DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_len[7:0]                       ), //i
    .io_input_ar_payload_size      (DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_size[2:0]                      ), //i
    .io_input_ar_payload_burst     (DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_burst[1:0]                     ), //i
    .io_input_ar_payload_prot      (DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_prot[2:0]                      ), //i
    .io_input_r_valid              (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_valid                  ), //o
    .io_input_r_ready              (DataCachePlugin_setup_dcacheMaster_readOnly_r_ready                                   ), //i
    .io_input_r_payload_data       (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_data[31:0]     ), //o
    .io_input_r_payload_id         (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_id[2:0]        ), //o
    .io_input_r_payload_resp       (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_resp[1:0]      ), //o
    .io_input_r_payload_last       (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_last           ), //o
    .io_outputs_0_ar_valid         (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_valid             ), //o
    .io_outputs_0_ar_ready         (io_outputs_0_ar_validPipe_fire_2                                                      ), //i
    .io_outputs_0_ar_payload_addr  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_addr[31:0]), //o
    .io_outputs_0_ar_payload_id    (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_id[2:0]   ), //o
    .io_outputs_0_ar_payload_len   (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_len[7:0]  ), //o
    .io_outputs_0_ar_payload_size  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_size[2:0] ), //o
    .io_outputs_0_ar_payload_burst (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_burst[1:0]), //o
    .io_outputs_0_ar_payload_prot  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_prot[2:0] ), //o
    .io_outputs_0_r_valid          (axi4ReadOnlyArbiter_3_io_inputs_2_r_valid                                             ), //i
    .io_outputs_0_r_ready          (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_r_ready              ), //o
    .io_outputs_0_r_payload_data   (axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_data[31:0]                                ), //i
    .io_outputs_0_r_payload_id     (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_r_payload_id[2:0]    ), //i
    .io_outputs_0_r_payload_resp   (axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_resp[1:0]                                 ), //i
    .io_outputs_0_r_payload_last   (axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_last                                      ), //i
    .io_outputs_1_ar_valid         (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_valid             ), //o
    .io_outputs_1_ar_ready         (io_outputs_1_ar_validPipe_fire_2                                                      ), //i
    .io_outputs_1_ar_payload_addr  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_addr[31:0]), //o
    .io_outputs_1_ar_payload_id    (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_id[2:0]   ), //o
    .io_outputs_1_ar_payload_len   (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_len[7:0]  ), //o
    .io_outputs_1_ar_payload_size  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_size[2:0] ), //o
    .io_outputs_1_ar_payload_burst (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_burst[1:0]), //o
    .io_outputs_1_ar_payload_prot  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_prot[2:0] ), //o
    .io_outputs_1_r_valid          (axi4ReadOnlyArbiter_4_io_inputs_2_r_valid                                             ), //i
    .io_outputs_1_r_ready          (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_r_ready              ), //o
    .io_outputs_1_r_payload_data   (axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_data[31:0]                                ), //i
    .io_outputs_1_r_payload_id     (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_r_payload_id[2:0]    ), //i
    .io_outputs_1_r_payload_resp   (axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_resp[1:0]                                 ), //i
    .io_outputs_1_r_payload_last   (axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_last                                      ), //i
    .io_outputs_2_ar_valid         (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_valid             ), //o
    .io_outputs_2_ar_ready         (io_outputs_2_ar_validPipe_fire_2                                                      ), //i
    .io_outputs_2_ar_payload_addr  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_addr[31:0]), //o
    .io_outputs_2_ar_payload_id    (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_id[2:0]   ), //o
    .io_outputs_2_ar_payload_len   (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_len[7:0]  ), //o
    .io_outputs_2_ar_payload_size  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_size[2:0] ), //o
    .io_outputs_2_ar_payload_burst (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_burst[1:0]), //o
    .io_outputs_2_ar_payload_prot  (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_prot[2:0] ), //o
    .io_outputs_2_r_valid          (axi4ReadOnlyArbiter_5_io_inputs_2_r_valid                                             ), //i
    .io_outputs_2_r_ready          (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_r_ready              ), //o
    .io_outputs_2_r_payload_data   (axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_data[31:0]                                ), //i
    .io_outputs_2_r_payload_id     (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_r_payload_id[2:0]    ), //i
    .io_outputs_2_r_payload_resp   (axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_resp[1:0]                                 ), //i
    .io_outputs_2_r_payload_last   (axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_last                                      ), //i
    .clk                           (clk                                                                                   ), //i
    .reset                         (reset                                                                                 )  //i
  );
  Axi4WriteOnlyDecoder_2 DataCachePlugin_setup_dcacheMaster_writeOnly_decoder (
    .io_input_aw_valid             (DataCachePlugin_setup_dcacheMaster_writeOnly_aw_valid                                  ), //i
    .io_input_aw_ready             (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_aw_ready                 ), //o
    .io_input_aw_payload_addr      (DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_addr[31:0]                     ), //i
    .io_input_aw_payload_id        (DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_id[2:0]                        ), //i
    .io_input_aw_payload_len       (DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_len[7:0]                       ), //i
    .io_input_aw_payload_size      (DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_size[2:0]                      ), //i
    .io_input_aw_payload_burst     (DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_burst[1:0]                     ), //i
    .io_input_aw_payload_prot      (DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_prot[2:0]                      ), //i
    .io_input_w_valid              (DataCachePlugin_setup_dcacheMaster_writeOnly_w_valid                                   ), //i
    .io_input_w_ready              (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_w_ready                  ), //o
    .io_input_w_payload_data       (DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_data[31:0]                      ), //i
    .io_input_w_payload_strb       (DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_strb[3:0]                       ), //i
    .io_input_w_payload_last       (DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_last                            ), //i
    .io_input_b_valid              (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_valid                  ), //o
    .io_input_b_ready              (DataCachePlugin_setup_dcacheMaster_writeOnly_b_ready                                   ), //i
    .io_input_b_payload_id         (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_payload_id[2:0]        ), //o
    .io_input_b_payload_resp       (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_payload_resp[1:0]      ), //o
    .io_outputs_0_aw_valid         (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_valid             ), //o
    .io_outputs_0_aw_ready         (io_outputs_0_aw_validPipe_fire_2                                                       ), //i
    .io_outputs_0_aw_payload_addr  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_addr[31:0]), //o
    .io_outputs_0_aw_payload_id    (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_id[2:0]   ), //o
    .io_outputs_0_aw_payload_len   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_len[7:0]  ), //o
    .io_outputs_0_aw_payload_size  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_size[2:0] ), //o
    .io_outputs_0_aw_payload_burst (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_burst[1:0]), //o
    .io_outputs_0_aw_payload_prot  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_prot[2:0] ), //o
    .io_outputs_0_w_valid          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_valid              ), //o
    .io_outputs_0_w_ready          (axi4WriteOnlyArbiter_3_io_inputs_2_w_ready                                             ), //i
    .io_outputs_0_w_payload_data   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_data[31:0] ), //o
    .io_outputs_0_w_payload_strb   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]  ), //o
    .io_outputs_0_w_payload_last   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_last       ), //o
    .io_outputs_0_b_valid          (axi4WriteOnlyArbiter_3_io_inputs_2_b_valid                                             ), //i
    .io_outputs_0_b_ready          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_b_ready              ), //o
    .io_outputs_0_b_payload_id     (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_b_payload_id[2:0]    ), //i
    .io_outputs_0_b_payload_resp   (axi4WriteOnlyArbiter_3_io_inputs_2_b_payload_resp[1:0]                                 ), //i
    .io_outputs_1_aw_valid         (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_valid             ), //o
    .io_outputs_1_aw_ready         (io_outputs_1_aw_validPipe_fire_2                                                       ), //i
    .io_outputs_1_aw_payload_addr  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_addr[31:0]), //o
    .io_outputs_1_aw_payload_id    (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_id[2:0]   ), //o
    .io_outputs_1_aw_payload_len   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_len[7:0]  ), //o
    .io_outputs_1_aw_payload_size  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_size[2:0] ), //o
    .io_outputs_1_aw_payload_burst (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_burst[1:0]), //o
    .io_outputs_1_aw_payload_prot  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_prot[2:0] ), //o
    .io_outputs_1_w_valid          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_valid              ), //o
    .io_outputs_1_w_ready          (axi4WriteOnlyArbiter_4_io_inputs_2_w_ready                                             ), //i
    .io_outputs_1_w_payload_data   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_data[31:0] ), //o
    .io_outputs_1_w_payload_strb   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_strb[3:0]  ), //o
    .io_outputs_1_w_payload_last   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_last       ), //o
    .io_outputs_1_b_valid          (axi4WriteOnlyArbiter_4_io_inputs_2_b_valid                                             ), //i
    .io_outputs_1_b_ready          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_b_ready              ), //o
    .io_outputs_1_b_payload_id     (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_b_payload_id[2:0]    ), //i
    .io_outputs_1_b_payload_resp   (axi4WriteOnlyArbiter_4_io_inputs_2_b_payload_resp[1:0]                                 ), //i
    .io_outputs_2_aw_valid         (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_valid             ), //o
    .io_outputs_2_aw_ready         (io_outputs_2_aw_validPipe_fire_2                                                       ), //i
    .io_outputs_2_aw_payload_addr  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_addr[31:0]), //o
    .io_outputs_2_aw_payload_id    (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_id[2:0]   ), //o
    .io_outputs_2_aw_payload_len   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_len[7:0]  ), //o
    .io_outputs_2_aw_payload_size  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_size[2:0] ), //o
    .io_outputs_2_aw_payload_burst (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_burst[1:0]), //o
    .io_outputs_2_aw_payload_prot  (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_prot[2:0] ), //o
    .io_outputs_2_w_valid          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_valid              ), //o
    .io_outputs_2_w_ready          (axi4WriteOnlyArbiter_5_io_inputs_2_w_ready                                             ), //i
    .io_outputs_2_w_payload_data   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_data[31:0] ), //o
    .io_outputs_2_w_payload_strb   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_strb[3:0]  ), //o
    .io_outputs_2_w_payload_last   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_last       ), //o
    .io_outputs_2_b_valid          (axi4WriteOnlyArbiter_5_io_inputs_2_b_valid                                             ), //i
    .io_outputs_2_b_ready          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_b_ready              ), //o
    .io_outputs_2_b_payload_id     (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_b_payload_id[2:0]    ), //i
    .io_outputs_2_b_payload_resp   (axi4WriteOnlyArbiter_5_io_inputs_2_b_payload_resp[1:0]                                 ), //i
    .clk                           (clk                                                                                    ), //i
    .reset                         (reset                                                                                  )  //i
  );
  Axi4ReadOnlyDecoder CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder (
    .io_input_ar_valid             (CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_valid                                  ), //i
    .io_input_ar_ready             (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_ar_ready                 ), //o
    .io_input_ar_payload_addr      (CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_addr[31:0]                     ), //i
    .io_input_ar_payload_id        (CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_id[3:0]                        ), //i
    .io_input_ar_payload_len       (CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_len[7:0]                       ), //i
    .io_input_ar_payload_size      (CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_size[2:0]                      ), //i
    .io_input_ar_payload_burst     (CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_burst[1:0]                     ), //i
    .io_input_r_valid              (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_valid                  ), //o
    .io_input_r_ready              (CoreMemSysPlugin_logic_roMasters_0_readOnly_r_ready                                   ), //i
    .io_input_r_payload_data       (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_data[31:0]     ), //o
    .io_input_r_payload_id         (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_id[3:0]        ), //o
    .io_input_r_payload_resp       (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_resp[1:0]      ), //o
    .io_input_r_payload_last       (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_last           ), //o
    .io_outputs_0_ar_valid         (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_valid             ), //o
    .io_outputs_0_ar_ready         (io_outputs_0_ar_validPipe_fire_3                                                      ), //i
    .io_outputs_0_ar_payload_addr  (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_addr[31:0]), //o
    .io_outputs_0_ar_payload_id    (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_id[3:0]   ), //o
    .io_outputs_0_ar_payload_len   (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_len[7:0]  ), //o
    .io_outputs_0_ar_payload_size  (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_size[2:0] ), //o
    .io_outputs_0_ar_payload_burst (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_burst[1:0]), //o
    .io_outputs_0_r_valid          (axi4ReadOnlyArbiter_3_io_inputs_3_r_valid                                             ), //i
    .io_outputs_0_r_ready          (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_r_ready              ), //o
    .io_outputs_0_r_payload_data   (axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_data[31:0]                                ), //i
    .io_outputs_0_r_payload_id     (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_r_payload_id[3:0]    ), //i
    .io_outputs_0_r_payload_resp   (axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_resp[1:0]                                 ), //i
    .io_outputs_0_r_payload_last   (axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_last                                      ), //i
    .io_outputs_1_ar_valid         (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_valid             ), //o
    .io_outputs_1_ar_ready         (io_outputs_1_ar_validPipe_fire_3                                                      ), //i
    .io_outputs_1_ar_payload_addr  (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_addr[31:0]), //o
    .io_outputs_1_ar_payload_id    (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_id[3:0]   ), //o
    .io_outputs_1_ar_payload_len   (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_len[7:0]  ), //o
    .io_outputs_1_ar_payload_size  (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_size[2:0] ), //o
    .io_outputs_1_ar_payload_burst (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_burst[1:0]), //o
    .io_outputs_1_r_valid          (axi4ReadOnlyArbiter_4_io_inputs_3_r_valid                                             ), //i
    .io_outputs_1_r_ready          (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_r_ready              ), //o
    .io_outputs_1_r_payload_data   (axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_data[31:0]                                ), //i
    .io_outputs_1_r_payload_id     (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_r_payload_id[3:0]    ), //i
    .io_outputs_1_r_payload_resp   (axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_resp[1:0]                                 ), //i
    .io_outputs_1_r_payload_last   (axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_last                                      ), //i
    .io_outputs_2_ar_valid         (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_valid             ), //o
    .io_outputs_2_ar_ready         (io_outputs_2_ar_validPipe_fire_3                                                      ), //i
    .io_outputs_2_ar_payload_addr  (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_addr[31:0]), //o
    .io_outputs_2_ar_payload_id    (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_id[3:0]   ), //o
    .io_outputs_2_ar_payload_len   (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_len[7:0]  ), //o
    .io_outputs_2_ar_payload_size  (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_size[2:0] ), //o
    .io_outputs_2_ar_payload_burst (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_burst[1:0]), //o
    .io_outputs_2_r_valid          (axi4ReadOnlyArbiter_5_io_inputs_3_r_valid                                             ), //i
    .io_outputs_2_r_ready          (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_r_ready              ), //o
    .io_outputs_2_r_payload_data   (axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_data[31:0]                                ), //i
    .io_outputs_2_r_payload_id     (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_r_payload_id[3:0]    ), //i
    .io_outputs_2_r_payload_resp   (axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_resp[1:0]                                 ), //i
    .io_outputs_2_r_payload_last   (axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_last                                      ), //i
    .clk                           (clk                                                                                   ), //i
    .reset                         (reset                                                                                 )  //i
  );
  Axi4WriteOnlyDecoder CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder (
    .io_input_aw_valid             (CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_valid                                  ), //i
    .io_input_aw_ready             (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_aw_ready                 ), //o
    .io_input_aw_payload_addr      (CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_addr[31:0]                     ), //i
    .io_input_aw_payload_id        (CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_id[3:0]                        ), //i
    .io_input_aw_payload_len       (CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_len[7:0]                       ), //i
    .io_input_aw_payload_size      (CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_size[2:0]                      ), //i
    .io_input_aw_payload_burst     (CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_burst[1:0]                     ), //i
    .io_input_w_valid              (CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_valid                                   ), //i
    .io_input_w_ready              (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_w_ready                  ), //o
    .io_input_w_payload_data       (CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_data[31:0]                      ), //i
    .io_input_w_payload_strb       (CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_strb[3:0]                       ), //i
    .io_input_w_payload_last       (CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_last                            ), //i
    .io_input_b_valid              (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_valid                  ), //o
    .io_input_b_ready              (CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_ready                                   ), //i
    .io_input_b_payload_id         (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_payload_id[3:0]        ), //o
    .io_input_b_payload_resp       (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_payload_resp[1:0]      ), //o
    .io_outputs_0_aw_valid         (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_valid             ), //o
    .io_outputs_0_aw_ready         (io_outputs_0_aw_validPipe_fire_3                                                       ), //i
    .io_outputs_0_aw_payload_addr  (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_addr[31:0]), //o
    .io_outputs_0_aw_payload_id    (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_id[3:0]   ), //o
    .io_outputs_0_aw_payload_len   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_len[7:0]  ), //o
    .io_outputs_0_aw_payload_size  (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_size[2:0] ), //o
    .io_outputs_0_aw_payload_burst (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_burst[1:0]), //o
    .io_outputs_0_w_valid          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_valid              ), //o
    .io_outputs_0_w_ready          (axi4WriteOnlyArbiter_3_io_inputs_3_w_ready                                             ), //i
    .io_outputs_0_w_payload_data   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_data[31:0] ), //o
    .io_outputs_0_w_payload_strb   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]  ), //o
    .io_outputs_0_w_payload_last   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_last       ), //o
    .io_outputs_0_b_valid          (axi4WriteOnlyArbiter_3_io_inputs_3_b_valid                                             ), //i
    .io_outputs_0_b_ready          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_b_ready              ), //o
    .io_outputs_0_b_payload_id     (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_b_payload_id[3:0]    ), //i
    .io_outputs_0_b_payload_resp   (axi4WriteOnlyArbiter_3_io_inputs_3_b_payload_resp[1:0]                                 ), //i
    .io_outputs_1_aw_valid         (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_valid             ), //o
    .io_outputs_1_aw_ready         (io_outputs_1_aw_validPipe_fire_3                                                       ), //i
    .io_outputs_1_aw_payload_addr  (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_addr[31:0]), //o
    .io_outputs_1_aw_payload_id    (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_id[3:0]   ), //o
    .io_outputs_1_aw_payload_len   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_len[7:0]  ), //o
    .io_outputs_1_aw_payload_size  (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_size[2:0] ), //o
    .io_outputs_1_aw_payload_burst (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_burst[1:0]), //o
    .io_outputs_1_w_valid          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_valid              ), //o
    .io_outputs_1_w_ready          (axi4WriteOnlyArbiter_4_io_inputs_3_w_ready                                             ), //i
    .io_outputs_1_w_payload_data   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_data[31:0] ), //o
    .io_outputs_1_w_payload_strb   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_strb[3:0]  ), //o
    .io_outputs_1_w_payload_last   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_last       ), //o
    .io_outputs_1_b_valid          (axi4WriteOnlyArbiter_4_io_inputs_3_b_valid                                             ), //i
    .io_outputs_1_b_ready          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_b_ready              ), //o
    .io_outputs_1_b_payload_id     (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_b_payload_id[3:0]    ), //i
    .io_outputs_1_b_payload_resp   (axi4WriteOnlyArbiter_4_io_inputs_3_b_payload_resp[1:0]                                 ), //i
    .io_outputs_2_aw_valid         (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_valid             ), //o
    .io_outputs_2_aw_ready         (io_outputs_2_aw_validPipe_fire_3                                                       ), //i
    .io_outputs_2_aw_payload_addr  (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_addr[31:0]), //o
    .io_outputs_2_aw_payload_id    (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_id[3:0]   ), //o
    .io_outputs_2_aw_payload_len   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_len[7:0]  ), //o
    .io_outputs_2_aw_payload_size  (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_size[2:0] ), //o
    .io_outputs_2_aw_payload_burst (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_burst[1:0]), //o
    .io_outputs_2_w_valid          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_valid              ), //o
    .io_outputs_2_w_ready          (axi4WriteOnlyArbiter_5_io_inputs_3_w_ready                                             ), //i
    .io_outputs_2_w_payload_data   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_data[31:0] ), //o
    .io_outputs_2_w_payload_strb   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_strb[3:0]  ), //o
    .io_outputs_2_w_payload_last   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_last       ), //o
    .io_outputs_2_b_valid          (axi4WriteOnlyArbiter_5_io_inputs_3_b_valid                                             ), //i
    .io_outputs_2_b_ready          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_b_ready              ), //o
    .io_outputs_2_b_payload_id     (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_b_payload_id[3:0]    ), //i
    .io_outputs_2_b_payload_resp   (axi4WriteOnlyArbiter_5_io_inputs_3_b_payload_resp[1:0]                                 ), //i
    .clk                           (clk                                                                                    ), //i
    .reset                         (reset                                                                                  )  //i
  );
  Axi4ReadOnlyArbiter axi4ReadOnlyArbiter_3 (
    .io_inputs_0_ar_valid         (io_outputs_0_ar_validPipe_valid                                         ), //i
    .io_inputs_0_ar_ready         (axi4ReadOnlyArbiter_3_io_inputs_0_ar_ready                              ), //o
    .io_inputs_0_ar_payload_addr  (io_outputs_0_ar_validPipe_payload_addr[31:0]                            ), //i
    .io_inputs_0_ar_payload_id    (axi4ReadOnlyArbiter_3_io_inputs_0_ar_payload_id[4:0]                    ), //i
    .io_inputs_0_ar_payload_len   (io_outputs_0_ar_validPipe_payload_len[7:0]                              ), //i
    .io_inputs_0_ar_payload_size  (io_outputs_0_ar_validPipe_payload_size[2:0]                             ), //i
    .io_inputs_0_ar_payload_burst (io_outputs_0_ar_validPipe_payload_burst[1:0]                            ), //i
    .io_inputs_0_r_valid          (axi4ReadOnlyArbiter_3_io_inputs_0_r_valid                               ), //o
    .io_inputs_0_r_ready          (io_axiOut_readOnly_decoder_io_outputs_0_r_ready                         ), //i
    .io_inputs_0_r_payload_data   (axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_data[31:0]                  ), //o
    .io_inputs_0_r_payload_id     (axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_id[4:0]                     ), //o
    .io_inputs_0_r_payload_resp   (axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_resp[1:0]                   ), //o
    .io_inputs_0_r_payload_last   (axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_last                        ), //o
    .io_inputs_1_ar_valid         (io_outputs_0_ar_validPipe_valid_1                                       ), //i
    .io_inputs_1_ar_ready         (axi4ReadOnlyArbiter_3_io_inputs_1_ar_ready                              ), //o
    .io_inputs_1_ar_payload_addr  (io_outputs_0_ar_validPipe_payload_addr_1[31:0]                          ), //i
    .io_inputs_1_ar_payload_id    (axi4ReadOnlyArbiter_3_io_inputs_1_ar_payload_id[4:0]                    ), //i
    .io_inputs_1_ar_payload_len   (io_outputs_0_ar_validPipe_payload_len_1[7:0]                            ), //i
    .io_inputs_1_ar_payload_size  (io_outputs_0_ar_validPipe_payload_size_1[2:0]                           ), //i
    .io_inputs_1_ar_payload_burst (io_outputs_0_ar_validPipe_payload_burst_1[1:0]                          ), //i
    .io_inputs_1_r_valid          (axi4ReadOnlyArbiter_3_io_inputs_1_r_valid                               ), //o
    .io_inputs_1_r_ready          (io_axiOut_readOnly_decoder_1_io_outputs_0_r_ready                       ), //i
    .io_inputs_1_r_payload_data   (axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_data[31:0]                  ), //o
    .io_inputs_1_r_payload_id     (axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_id[4:0]                     ), //o
    .io_inputs_1_r_payload_resp   (axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_resp[1:0]                   ), //o
    .io_inputs_1_r_payload_last   (axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_last                        ), //o
    .io_inputs_2_ar_valid         (io_outputs_0_ar_validPipe_valid_2                                       ), //i
    .io_inputs_2_ar_ready         (axi4ReadOnlyArbiter_3_io_inputs_2_ar_ready                              ), //o
    .io_inputs_2_ar_payload_addr  (io_outputs_0_ar_validPipe_payload_addr_2[31:0]                          ), //i
    .io_inputs_2_ar_payload_id    (axi4ReadOnlyArbiter_3_io_inputs_2_ar_payload_id[4:0]                    ), //i
    .io_inputs_2_ar_payload_len   (io_outputs_0_ar_validPipe_payload_len_2[7:0]                            ), //i
    .io_inputs_2_ar_payload_size  (io_outputs_0_ar_validPipe_payload_size_2[2:0]                           ), //i
    .io_inputs_2_ar_payload_burst (io_outputs_0_ar_validPipe_payload_burst_2[1:0]                          ), //i
    .io_inputs_2_r_valid          (axi4ReadOnlyArbiter_3_io_inputs_2_r_valid                               ), //o
    .io_inputs_2_r_ready          (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_r_ready), //i
    .io_inputs_2_r_payload_data   (axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_data[31:0]                  ), //o
    .io_inputs_2_r_payload_id     (axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_id[4:0]                     ), //o
    .io_inputs_2_r_payload_resp   (axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_resp[1:0]                   ), //o
    .io_inputs_2_r_payload_last   (axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_last                        ), //o
    .io_inputs_3_ar_valid         (io_outputs_0_ar_validPipe_valid_3                                       ), //i
    .io_inputs_3_ar_ready         (axi4ReadOnlyArbiter_3_io_inputs_3_ar_ready                              ), //o
    .io_inputs_3_ar_payload_addr  (io_outputs_0_ar_validPipe_payload_addr_3[31:0]                          ), //i
    .io_inputs_3_ar_payload_id    (axi4ReadOnlyArbiter_3_io_inputs_3_ar_payload_id[4:0]                    ), //i
    .io_inputs_3_ar_payload_len   (io_outputs_0_ar_validPipe_payload_len_3[7:0]                            ), //i
    .io_inputs_3_ar_payload_size  (io_outputs_0_ar_validPipe_payload_size_3[2:0]                           ), //i
    .io_inputs_3_ar_payload_burst (io_outputs_0_ar_validPipe_payload_burst_3[1:0]                          ), //i
    .io_inputs_3_r_valid          (axi4ReadOnlyArbiter_3_io_inputs_3_r_valid                               ), //o
    .io_inputs_3_r_ready          (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_r_ready), //i
    .io_inputs_3_r_payload_data   (axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_data[31:0]                  ), //o
    .io_inputs_3_r_payload_id     (axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_id[4:0]                     ), //o
    .io_inputs_3_r_payload_resp   (axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_resp[1:0]                   ), //o
    .io_inputs_3_r_payload_last   (axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_last                        ), //o
    .io_output_ar_valid           (axi4ReadOnlyArbiter_3_io_output_ar_valid                                ), //o
    .io_output_ar_ready           (CoreMemSysPlugin_hw_baseramCtrl_io_axi_ar_ready                         ), //i
    .io_output_ar_payload_addr    (axi4ReadOnlyArbiter_3_io_output_ar_payload_addr[31:0]                   ), //o
    .io_output_ar_payload_id      (axi4ReadOnlyArbiter_3_io_output_ar_payload_id[6:0]                      ), //o
    .io_output_ar_payload_len     (axi4ReadOnlyArbiter_3_io_output_ar_payload_len[7:0]                     ), //o
    .io_output_ar_payload_size    (axi4ReadOnlyArbiter_3_io_output_ar_payload_size[2:0]                    ), //o
    .io_output_ar_payload_burst   (axi4ReadOnlyArbiter_3_io_output_ar_payload_burst[1:0]                   ), //o
    .io_output_r_valid            (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_valid                          ), //i
    .io_output_r_ready            (axi4ReadOnlyArbiter_3_io_output_r_ready                                 ), //o
    .io_output_r_payload_data     (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_data[31:0]             ), //i
    .io_output_r_payload_id       (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_id[6:0]                ), //i
    .io_output_r_payload_resp     (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_resp[1:0]              ), //i
    .io_output_r_payload_last     (CoreMemSysPlugin_hw_baseramCtrl_io_axi_r_payload_last                   ), //i
    .clk                          (clk                                                                     ), //i
    .reset                        (reset                                                                   )  //i
  );
  Axi4WriteOnlyArbiter axi4WriteOnlyArbiter_3 (
    .io_inputs_0_aw_valid         (io_outputs_0_aw_validPipe_valid                                                       ), //i
    .io_inputs_0_aw_ready         (axi4WriteOnlyArbiter_3_io_inputs_0_aw_ready                                           ), //o
    .io_inputs_0_aw_payload_addr  (io_outputs_0_aw_validPipe_payload_addr[31:0]                                          ), //i
    .io_inputs_0_aw_payload_id    (axi4WriteOnlyArbiter_3_io_inputs_0_aw_payload_id[4:0]                                 ), //i
    .io_inputs_0_aw_payload_len   (io_outputs_0_aw_validPipe_payload_len[7:0]                                            ), //i
    .io_inputs_0_aw_payload_size  (io_outputs_0_aw_validPipe_payload_size[2:0]                                           ), //i
    .io_inputs_0_aw_payload_burst (io_outputs_0_aw_validPipe_payload_burst[1:0]                                          ), //i
    .io_inputs_0_w_valid          (io_axiOut_writeOnly_decoder_io_outputs_0_w_valid                                      ), //i
    .io_inputs_0_w_ready          (axi4WriteOnlyArbiter_3_io_inputs_0_w_ready                                            ), //o
    .io_inputs_0_w_payload_data   (io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]                         ), //i
    .io_inputs_0_w_payload_strb   (io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]                          ), //i
    .io_inputs_0_w_payload_last   (io_axiOut_writeOnly_decoder_io_outputs_0_w_payload_last                               ), //i
    .io_inputs_0_b_valid          (axi4WriteOnlyArbiter_3_io_inputs_0_b_valid                                            ), //o
    .io_inputs_0_b_ready          (io_axiOut_writeOnly_decoder_io_outputs_0_b_ready                                      ), //i
    .io_inputs_0_b_payload_id     (axi4WriteOnlyArbiter_3_io_inputs_0_b_payload_id[4:0]                                  ), //o
    .io_inputs_0_b_payload_resp   (axi4WriteOnlyArbiter_3_io_inputs_0_b_payload_resp[1:0]                                ), //o
    .io_inputs_1_aw_valid         (io_outputs_0_aw_validPipe_valid_1                                                     ), //i
    .io_inputs_1_aw_ready         (axi4WriteOnlyArbiter_3_io_inputs_1_aw_ready                                           ), //o
    .io_inputs_1_aw_payload_addr  (io_outputs_0_aw_validPipe_payload_addr_1[31:0]                                        ), //i
    .io_inputs_1_aw_payload_id    (axi4WriteOnlyArbiter_3_io_inputs_1_aw_payload_id[4:0]                                 ), //i
    .io_inputs_1_aw_payload_len   (io_outputs_0_aw_validPipe_payload_len_1[7:0]                                          ), //i
    .io_inputs_1_aw_payload_size  (io_outputs_0_aw_validPipe_payload_size_1[2:0]                                         ), //i
    .io_inputs_1_aw_payload_burst (io_outputs_0_aw_validPipe_payload_burst_1[1:0]                                        ), //i
    .io_inputs_1_w_valid          (io_axiOut_writeOnly_decoder_1_io_outputs_0_w_valid                                    ), //i
    .io_inputs_1_w_ready          (axi4WriteOnlyArbiter_3_io_inputs_1_w_ready                                            ), //o
    .io_inputs_1_w_payload_data   (io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_data[31:0]                       ), //i
    .io_inputs_1_w_payload_strb   (io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_strb[3:0]                        ), //i
    .io_inputs_1_w_payload_last   (io_axiOut_writeOnly_decoder_1_io_outputs_0_w_payload_last                             ), //i
    .io_inputs_1_b_valid          (axi4WriteOnlyArbiter_3_io_inputs_1_b_valid                                            ), //o
    .io_inputs_1_b_ready          (io_axiOut_writeOnly_decoder_1_io_outputs_0_b_ready                                    ), //i
    .io_inputs_1_b_payload_id     (axi4WriteOnlyArbiter_3_io_inputs_1_b_payload_id[4:0]                                  ), //o
    .io_inputs_1_b_payload_resp   (axi4WriteOnlyArbiter_3_io_inputs_1_b_payload_resp[1:0]                                ), //o
    .io_inputs_2_aw_valid         (io_outputs_0_aw_validPipe_valid_2                                                     ), //i
    .io_inputs_2_aw_ready         (axi4WriteOnlyArbiter_3_io_inputs_2_aw_ready                                           ), //o
    .io_inputs_2_aw_payload_addr  (io_outputs_0_aw_validPipe_payload_addr_2[31:0]                                        ), //i
    .io_inputs_2_aw_payload_id    (axi4WriteOnlyArbiter_3_io_inputs_2_aw_payload_id[4:0]                                 ), //i
    .io_inputs_2_aw_payload_len   (io_outputs_0_aw_validPipe_payload_len_2[7:0]                                          ), //i
    .io_inputs_2_aw_payload_size  (io_outputs_0_aw_validPipe_payload_size_2[2:0]                                         ), //i
    .io_inputs_2_aw_payload_burst (io_outputs_0_aw_validPipe_payload_burst_2[1:0]                                        ), //i
    .io_inputs_2_w_valid          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_valid             ), //i
    .io_inputs_2_w_ready          (axi4WriteOnlyArbiter_3_io_inputs_2_w_ready                                            ), //o
    .io_inputs_2_w_payload_data   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]), //i
    .io_inputs_2_w_payload_strb   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0] ), //i
    .io_inputs_2_w_payload_last   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_w_payload_last      ), //i
    .io_inputs_2_b_valid          (axi4WriteOnlyArbiter_3_io_inputs_2_b_valid                                            ), //o
    .io_inputs_2_b_ready          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_b_ready             ), //i
    .io_inputs_2_b_payload_id     (axi4WriteOnlyArbiter_3_io_inputs_2_b_payload_id[4:0]                                  ), //o
    .io_inputs_2_b_payload_resp   (axi4WriteOnlyArbiter_3_io_inputs_2_b_payload_resp[1:0]                                ), //o
    .io_inputs_3_aw_valid         (io_outputs_0_aw_validPipe_valid_3                                                     ), //i
    .io_inputs_3_aw_ready         (axi4WriteOnlyArbiter_3_io_inputs_3_aw_ready                                           ), //o
    .io_inputs_3_aw_payload_addr  (io_outputs_0_aw_validPipe_payload_addr_3[31:0]                                        ), //i
    .io_inputs_3_aw_payload_id    (axi4WriteOnlyArbiter_3_io_inputs_3_aw_payload_id[4:0]                                 ), //i
    .io_inputs_3_aw_payload_len   (io_outputs_0_aw_validPipe_payload_len_3[7:0]                                          ), //i
    .io_inputs_3_aw_payload_size  (io_outputs_0_aw_validPipe_payload_size_3[2:0]                                         ), //i
    .io_inputs_3_aw_payload_burst (io_outputs_0_aw_validPipe_payload_burst_3[1:0]                                        ), //i
    .io_inputs_3_w_valid          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_valid             ), //i
    .io_inputs_3_w_ready          (axi4WriteOnlyArbiter_3_io_inputs_3_w_ready                                            ), //o
    .io_inputs_3_w_payload_data   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]), //i
    .io_inputs_3_w_payload_strb   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0] ), //i
    .io_inputs_3_w_payload_last   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_w_payload_last      ), //i
    .io_inputs_3_b_valid          (axi4WriteOnlyArbiter_3_io_inputs_3_b_valid                                            ), //o
    .io_inputs_3_b_ready          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_b_ready             ), //i
    .io_inputs_3_b_payload_id     (axi4WriteOnlyArbiter_3_io_inputs_3_b_payload_id[4:0]                                  ), //o
    .io_inputs_3_b_payload_resp   (axi4WriteOnlyArbiter_3_io_inputs_3_b_payload_resp[1:0]                                ), //o
    .io_output_aw_valid           (axi4WriteOnlyArbiter_3_io_output_aw_valid                                             ), //o
    .io_output_aw_ready           (CoreMemSysPlugin_hw_baseramCtrl_io_axi_aw_ready                                       ), //i
    .io_output_aw_payload_addr    (axi4WriteOnlyArbiter_3_io_output_aw_payload_addr[31:0]                                ), //o
    .io_output_aw_payload_id      (axi4WriteOnlyArbiter_3_io_output_aw_payload_id[6:0]                                   ), //o
    .io_output_aw_payload_len     (axi4WriteOnlyArbiter_3_io_output_aw_payload_len[7:0]                                  ), //o
    .io_output_aw_payload_size    (axi4WriteOnlyArbiter_3_io_output_aw_payload_size[2:0]                                 ), //o
    .io_output_aw_payload_burst   (axi4WriteOnlyArbiter_3_io_output_aw_payload_burst[1:0]                                ), //o
    .io_output_w_valid            (axi4WriteOnlyArbiter_3_io_output_w_valid                                              ), //o
    .io_output_w_ready            (CoreMemSysPlugin_hw_baseramCtrl_io_axi_w_ready                                        ), //i
    .io_output_w_payload_data     (axi4WriteOnlyArbiter_3_io_output_w_payload_data[31:0]                                 ), //o
    .io_output_w_payload_strb     (axi4WriteOnlyArbiter_3_io_output_w_payload_strb[3:0]                                  ), //o
    .io_output_w_payload_last     (axi4WriteOnlyArbiter_3_io_output_w_payload_last                                       ), //o
    .io_output_b_valid            (CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_valid                                        ), //i
    .io_output_b_ready            (axi4WriteOnlyArbiter_3_io_output_b_ready                                              ), //o
    .io_output_b_payload_id       (CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_payload_id[6:0]                              ), //i
    .io_output_b_payload_resp     (CoreMemSysPlugin_hw_baseramCtrl_io_axi_b_payload_resp[1:0]                            ), //i
    .clk                          (clk                                                                                   ), //i
    .reset                        (reset                                                                                 )  //i
  );
  Axi4ReadOnlyArbiter axi4ReadOnlyArbiter_4 (
    .io_inputs_0_ar_valid         (io_outputs_1_ar_validPipe_valid                                         ), //i
    .io_inputs_0_ar_ready         (axi4ReadOnlyArbiter_4_io_inputs_0_ar_ready                              ), //o
    .io_inputs_0_ar_payload_addr  (io_outputs_1_ar_validPipe_payload_addr[31:0]                            ), //i
    .io_inputs_0_ar_payload_id    (axi4ReadOnlyArbiter_4_io_inputs_0_ar_payload_id[4:0]                    ), //i
    .io_inputs_0_ar_payload_len   (io_outputs_1_ar_validPipe_payload_len[7:0]                              ), //i
    .io_inputs_0_ar_payload_size  (io_outputs_1_ar_validPipe_payload_size[2:0]                             ), //i
    .io_inputs_0_ar_payload_burst (io_outputs_1_ar_validPipe_payload_burst[1:0]                            ), //i
    .io_inputs_0_r_valid          (axi4ReadOnlyArbiter_4_io_inputs_0_r_valid                               ), //o
    .io_inputs_0_r_ready          (io_axiOut_readOnly_decoder_io_outputs_1_r_ready                         ), //i
    .io_inputs_0_r_payload_data   (axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_data[31:0]                  ), //o
    .io_inputs_0_r_payload_id     (axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_id[4:0]                     ), //o
    .io_inputs_0_r_payload_resp   (axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_resp[1:0]                   ), //o
    .io_inputs_0_r_payload_last   (axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_last                        ), //o
    .io_inputs_1_ar_valid         (io_outputs_1_ar_validPipe_valid_1                                       ), //i
    .io_inputs_1_ar_ready         (axi4ReadOnlyArbiter_4_io_inputs_1_ar_ready                              ), //o
    .io_inputs_1_ar_payload_addr  (io_outputs_1_ar_validPipe_payload_addr_1[31:0]                          ), //i
    .io_inputs_1_ar_payload_id    (axi4ReadOnlyArbiter_4_io_inputs_1_ar_payload_id[4:0]                    ), //i
    .io_inputs_1_ar_payload_len   (io_outputs_1_ar_validPipe_payload_len_1[7:0]                            ), //i
    .io_inputs_1_ar_payload_size  (io_outputs_1_ar_validPipe_payload_size_1[2:0]                           ), //i
    .io_inputs_1_ar_payload_burst (io_outputs_1_ar_validPipe_payload_burst_1[1:0]                          ), //i
    .io_inputs_1_r_valid          (axi4ReadOnlyArbiter_4_io_inputs_1_r_valid                               ), //o
    .io_inputs_1_r_ready          (io_axiOut_readOnly_decoder_1_io_outputs_1_r_ready                       ), //i
    .io_inputs_1_r_payload_data   (axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_data[31:0]                  ), //o
    .io_inputs_1_r_payload_id     (axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_id[4:0]                     ), //o
    .io_inputs_1_r_payload_resp   (axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_resp[1:0]                   ), //o
    .io_inputs_1_r_payload_last   (axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_last                        ), //o
    .io_inputs_2_ar_valid         (io_outputs_1_ar_validPipe_valid_2                                       ), //i
    .io_inputs_2_ar_ready         (axi4ReadOnlyArbiter_4_io_inputs_2_ar_ready                              ), //o
    .io_inputs_2_ar_payload_addr  (io_outputs_1_ar_validPipe_payload_addr_2[31:0]                          ), //i
    .io_inputs_2_ar_payload_id    (axi4ReadOnlyArbiter_4_io_inputs_2_ar_payload_id[4:0]                    ), //i
    .io_inputs_2_ar_payload_len   (io_outputs_1_ar_validPipe_payload_len_2[7:0]                            ), //i
    .io_inputs_2_ar_payload_size  (io_outputs_1_ar_validPipe_payload_size_2[2:0]                           ), //i
    .io_inputs_2_ar_payload_burst (io_outputs_1_ar_validPipe_payload_burst_2[1:0]                          ), //i
    .io_inputs_2_r_valid          (axi4ReadOnlyArbiter_4_io_inputs_2_r_valid                               ), //o
    .io_inputs_2_r_ready          (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_r_ready), //i
    .io_inputs_2_r_payload_data   (axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_data[31:0]                  ), //o
    .io_inputs_2_r_payload_id     (axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_id[4:0]                     ), //o
    .io_inputs_2_r_payload_resp   (axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_resp[1:0]                   ), //o
    .io_inputs_2_r_payload_last   (axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_last                        ), //o
    .io_inputs_3_ar_valid         (io_outputs_1_ar_validPipe_valid_3                                       ), //i
    .io_inputs_3_ar_ready         (axi4ReadOnlyArbiter_4_io_inputs_3_ar_ready                              ), //o
    .io_inputs_3_ar_payload_addr  (io_outputs_1_ar_validPipe_payload_addr_3[31:0]                          ), //i
    .io_inputs_3_ar_payload_id    (axi4ReadOnlyArbiter_4_io_inputs_3_ar_payload_id[4:0]                    ), //i
    .io_inputs_3_ar_payload_len   (io_outputs_1_ar_validPipe_payload_len_3[7:0]                            ), //i
    .io_inputs_3_ar_payload_size  (io_outputs_1_ar_validPipe_payload_size_3[2:0]                           ), //i
    .io_inputs_3_ar_payload_burst (io_outputs_1_ar_validPipe_payload_burst_3[1:0]                          ), //i
    .io_inputs_3_r_valid          (axi4ReadOnlyArbiter_4_io_inputs_3_r_valid                               ), //o
    .io_inputs_3_r_ready          (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_r_ready), //i
    .io_inputs_3_r_payload_data   (axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_data[31:0]                  ), //o
    .io_inputs_3_r_payload_id     (axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_id[4:0]                     ), //o
    .io_inputs_3_r_payload_resp   (axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_resp[1:0]                   ), //o
    .io_inputs_3_r_payload_last   (axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_last                        ), //o
    .io_output_ar_valid           (axi4ReadOnlyArbiter_4_io_output_ar_valid                                ), //o
    .io_output_ar_ready           (CoreMemSysPlugin_hw_extramCtrl_io_axi_ar_ready                          ), //i
    .io_output_ar_payload_addr    (axi4ReadOnlyArbiter_4_io_output_ar_payload_addr[31:0]                   ), //o
    .io_output_ar_payload_id      (axi4ReadOnlyArbiter_4_io_output_ar_payload_id[6:0]                      ), //o
    .io_output_ar_payload_len     (axi4ReadOnlyArbiter_4_io_output_ar_payload_len[7:0]                     ), //o
    .io_output_ar_payload_size    (axi4ReadOnlyArbiter_4_io_output_ar_payload_size[2:0]                    ), //o
    .io_output_ar_payload_burst   (axi4ReadOnlyArbiter_4_io_output_ar_payload_burst[1:0]                   ), //o
    .io_output_r_valid            (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_valid                           ), //i
    .io_output_r_ready            (axi4ReadOnlyArbiter_4_io_output_r_ready                                 ), //o
    .io_output_r_payload_data     (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_data[31:0]              ), //i
    .io_output_r_payload_id       (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_id[6:0]                 ), //i
    .io_output_r_payload_resp     (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_resp[1:0]               ), //i
    .io_output_r_payload_last     (CoreMemSysPlugin_hw_extramCtrl_io_axi_r_payload_last                    ), //i
    .clk                          (clk                                                                     ), //i
    .reset                        (reset                                                                   )  //i
  );
  Axi4WriteOnlyArbiter axi4WriteOnlyArbiter_4 (
    .io_inputs_0_aw_valid         (io_outputs_1_aw_validPipe_valid                                                       ), //i
    .io_inputs_0_aw_ready         (axi4WriteOnlyArbiter_4_io_inputs_0_aw_ready                                           ), //o
    .io_inputs_0_aw_payload_addr  (io_outputs_1_aw_validPipe_payload_addr[31:0]                                          ), //i
    .io_inputs_0_aw_payload_id    (axi4WriteOnlyArbiter_4_io_inputs_0_aw_payload_id[4:0]                                 ), //i
    .io_inputs_0_aw_payload_len   (io_outputs_1_aw_validPipe_payload_len[7:0]                                            ), //i
    .io_inputs_0_aw_payload_size  (io_outputs_1_aw_validPipe_payload_size[2:0]                                           ), //i
    .io_inputs_0_aw_payload_burst (io_outputs_1_aw_validPipe_payload_burst[1:0]                                          ), //i
    .io_inputs_0_w_valid          (io_axiOut_writeOnly_decoder_io_outputs_1_w_valid                                      ), //i
    .io_inputs_0_w_ready          (axi4WriteOnlyArbiter_4_io_inputs_0_w_ready                                            ), //o
    .io_inputs_0_w_payload_data   (io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_data[31:0]                         ), //i
    .io_inputs_0_w_payload_strb   (io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_strb[3:0]                          ), //i
    .io_inputs_0_w_payload_last   (io_axiOut_writeOnly_decoder_io_outputs_1_w_payload_last                               ), //i
    .io_inputs_0_b_valid          (axi4WriteOnlyArbiter_4_io_inputs_0_b_valid                                            ), //o
    .io_inputs_0_b_ready          (io_axiOut_writeOnly_decoder_io_outputs_1_b_ready                                      ), //i
    .io_inputs_0_b_payload_id     (axi4WriteOnlyArbiter_4_io_inputs_0_b_payload_id[4:0]                                  ), //o
    .io_inputs_0_b_payload_resp   (axi4WriteOnlyArbiter_4_io_inputs_0_b_payload_resp[1:0]                                ), //o
    .io_inputs_1_aw_valid         (io_outputs_1_aw_validPipe_valid_1                                                     ), //i
    .io_inputs_1_aw_ready         (axi4WriteOnlyArbiter_4_io_inputs_1_aw_ready                                           ), //o
    .io_inputs_1_aw_payload_addr  (io_outputs_1_aw_validPipe_payload_addr_1[31:0]                                        ), //i
    .io_inputs_1_aw_payload_id    (axi4WriteOnlyArbiter_4_io_inputs_1_aw_payload_id[4:0]                                 ), //i
    .io_inputs_1_aw_payload_len   (io_outputs_1_aw_validPipe_payload_len_1[7:0]                                          ), //i
    .io_inputs_1_aw_payload_size  (io_outputs_1_aw_validPipe_payload_size_1[2:0]                                         ), //i
    .io_inputs_1_aw_payload_burst (io_outputs_1_aw_validPipe_payload_burst_1[1:0]                                        ), //i
    .io_inputs_1_w_valid          (io_axiOut_writeOnly_decoder_1_io_outputs_1_w_valid                                    ), //i
    .io_inputs_1_w_ready          (axi4WriteOnlyArbiter_4_io_inputs_1_w_ready                                            ), //o
    .io_inputs_1_w_payload_data   (io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_data[31:0]                       ), //i
    .io_inputs_1_w_payload_strb   (io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_strb[3:0]                        ), //i
    .io_inputs_1_w_payload_last   (io_axiOut_writeOnly_decoder_1_io_outputs_1_w_payload_last                             ), //i
    .io_inputs_1_b_valid          (axi4WriteOnlyArbiter_4_io_inputs_1_b_valid                                            ), //o
    .io_inputs_1_b_ready          (io_axiOut_writeOnly_decoder_1_io_outputs_1_b_ready                                    ), //i
    .io_inputs_1_b_payload_id     (axi4WriteOnlyArbiter_4_io_inputs_1_b_payload_id[4:0]                                  ), //o
    .io_inputs_1_b_payload_resp   (axi4WriteOnlyArbiter_4_io_inputs_1_b_payload_resp[1:0]                                ), //o
    .io_inputs_2_aw_valid         (io_outputs_1_aw_validPipe_valid_2                                                     ), //i
    .io_inputs_2_aw_ready         (axi4WriteOnlyArbiter_4_io_inputs_2_aw_ready                                           ), //o
    .io_inputs_2_aw_payload_addr  (io_outputs_1_aw_validPipe_payload_addr_2[31:0]                                        ), //i
    .io_inputs_2_aw_payload_id    (axi4WriteOnlyArbiter_4_io_inputs_2_aw_payload_id[4:0]                                 ), //i
    .io_inputs_2_aw_payload_len   (io_outputs_1_aw_validPipe_payload_len_2[7:0]                                          ), //i
    .io_inputs_2_aw_payload_size  (io_outputs_1_aw_validPipe_payload_size_2[2:0]                                         ), //i
    .io_inputs_2_aw_payload_burst (io_outputs_1_aw_validPipe_payload_burst_2[1:0]                                        ), //i
    .io_inputs_2_w_valid          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_valid             ), //i
    .io_inputs_2_w_ready          (axi4WriteOnlyArbiter_4_io_inputs_2_w_ready                                            ), //o
    .io_inputs_2_w_payload_data   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_data[31:0]), //i
    .io_inputs_2_w_payload_strb   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_strb[3:0] ), //i
    .io_inputs_2_w_payload_last   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_w_payload_last      ), //i
    .io_inputs_2_b_valid          (axi4WriteOnlyArbiter_4_io_inputs_2_b_valid                                            ), //o
    .io_inputs_2_b_ready          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_b_ready             ), //i
    .io_inputs_2_b_payload_id     (axi4WriteOnlyArbiter_4_io_inputs_2_b_payload_id[4:0]                                  ), //o
    .io_inputs_2_b_payload_resp   (axi4WriteOnlyArbiter_4_io_inputs_2_b_payload_resp[1:0]                                ), //o
    .io_inputs_3_aw_valid         (io_outputs_1_aw_validPipe_valid_3                                                     ), //i
    .io_inputs_3_aw_ready         (axi4WriteOnlyArbiter_4_io_inputs_3_aw_ready                                           ), //o
    .io_inputs_3_aw_payload_addr  (io_outputs_1_aw_validPipe_payload_addr_3[31:0]                                        ), //i
    .io_inputs_3_aw_payload_id    (axi4WriteOnlyArbiter_4_io_inputs_3_aw_payload_id[4:0]                                 ), //i
    .io_inputs_3_aw_payload_len   (io_outputs_1_aw_validPipe_payload_len_3[7:0]                                          ), //i
    .io_inputs_3_aw_payload_size  (io_outputs_1_aw_validPipe_payload_size_3[2:0]                                         ), //i
    .io_inputs_3_aw_payload_burst (io_outputs_1_aw_validPipe_payload_burst_3[1:0]                                        ), //i
    .io_inputs_3_w_valid          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_valid             ), //i
    .io_inputs_3_w_ready          (axi4WriteOnlyArbiter_4_io_inputs_3_w_ready                                            ), //o
    .io_inputs_3_w_payload_data   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_data[31:0]), //i
    .io_inputs_3_w_payload_strb   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_strb[3:0] ), //i
    .io_inputs_3_w_payload_last   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_w_payload_last      ), //i
    .io_inputs_3_b_valid          (axi4WriteOnlyArbiter_4_io_inputs_3_b_valid                                            ), //o
    .io_inputs_3_b_ready          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_b_ready             ), //i
    .io_inputs_3_b_payload_id     (axi4WriteOnlyArbiter_4_io_inputs_3_b_payload_id[4:0]                                  ), //o
    .io_inputs_3_b_payload_resp   (axi4WriteOnlyArbiter_4_io_inputs_3_b_payload_resp[1:0]                                ), //o
    .io_output_aw_valid           (axi4WriteOnlyArbiter_4_io_output_aw_valid                                             ), //o
    .io_output_aw_ready           (CoreMemSysPlugin_hw_extramCtrl_io_axi_aw_ready                                        ), //i
    .io_output_aw_payload_addr    (axi4WriteOnlyArbiter_4_io_output_aw_payload_addr[31:0]                                ), //o
    .io_output_aw_payload_id      (axi4WriteOnlyArbiter_4_io_output_aw_payload_id[6:0]                                   ), //o
    .io_output_aw_payload_len     (axi4WriteOnlyArbiter_4_io_output_aw_payload_len[7:0]                                  ), //o
    .io_output_aw_payload_size    (axi4WriteOnlyArbiter_4_io_output_aw_payload_size[2:0]                                 ), //o
    .io_output_aw_payload_burst   (axi4WriteOnlyArbiter_4_io_output_aw_payload_burst[1:0]                                ), //o
    .io_output_w_valid            (axi4WriteOnlyArbiter_4_io_output_w_valid                                              ), //o
    .io_output_w_ready            (CoreMemSysPlugin_hw_extramCtrl_io_axi_w_ready                                         ), //i
    .io_output_w_payload_data     (axi4WriteOnlyArbiter_4_io_output_w_payload_data[31:0]                                 ), //o
    .io_output_w_payload_strb     (axi4WriteOnlyArbiter_4_io_output_w_payload_strb[3:0]                                  ), //o
    .io_output_w_payload_last     (axi4WriteOnlyArbiter_4_io_output_w_payload_last                                       ), //o
    .io_output_b_valid            (CoreMemSysPlugin_hw_extramCtrl_io_axi_b_valid                                         ), //i
    .io_output_b_ready            (axi4WriteOnlyArbiter_4_io_output_b_ready                                              ), //o
    .io_output_b_payload_id       (CoreMemSysPlugin_hw_extramCtrl_io_axi_b_payload_id[6:0]                               ), //i
    .io_output_b_payload_resp     (CoreMemSysPlugin_hw_extramCtrl_io_axi_b_payload_resp[1:0]                             ), //i
    .clk                          (clk                                                                                   ), //i
    .reset                        (reset                                                                                 )  //i
  );
  Axi4ReadOnlyArbiter axi4ReadOnlyArbiter_5 (
    .io_inputs_0_ar_valid         (io_outputs_2_ar_validPipe_valid                                         ), //i
    .io_inputs_0_ar_ready         (axi4ReadOnlyArbiter_5_io_inputs_0_ar_ready                              ), //o
    .io_inputs_0_ar_payload_addr  (io_outputs_2_ar_validPipe_payload_addr[31:0]                            ), //i
    .io_inputs_0_ar_payload_id    (axi4ReadOnlyArbiter_5_io_inputs_0_ar_payload_id[4:0]                    ), //i
    .io_inputs_0_ar_payload_len   (io_outputs_2_ar_validPipe_payload_len[7:0]                              ), //i
    .io_inputs_0_ar_payload_size  (io_outputs_2_ar_validPipe_payload_size[2:0]                             ), //i
    .io_inputs_0_ar_payload_burst (io_outputs_2_ar_validPipe_payload_burst[1:0]                            ), //i
    .io_inputs_0_r_valid          (axi4ReadOnlyArbiter_5_io_inputs_0_r_valid                               ), //o
    .io_inputs_0_r_ready          (io_axiOut_readOnly_decoder_io_outputs_2_r_ready                         ), //i
    .io_inputs_0_r_payload_data   (axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_data[31:0]                  ), //o
    .io_inputs_0_r_payload_id     (axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_id[4:0]                     ), //o
    .io_inputs_0_r_payload_resp   (axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_resp[1:0]                   ), //o
    .io_inputs_0_r_payload_last   (axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_last                        ), //o
    .io_inputs_1_ar_valid         (io_outputs_2_ar_validPipe_valid_1                                       ), //i
    .io_inputs_1_ar_ready         (axi4ReadOnlyArbiter_5_io_inputs_1_ar_ready                              ), //o
    .io_inputs_1_ar_payload_addr  (io_outputs_2_ar_validPipe_payload_addr_1[31:0]                          ), //i
    .io_inputs_1_ar_payload_id    (axi4ReadOnlyArbiter_5_io_inputs_1_ar_payload_id[4:0]                    ), //i
    .io_inputs_1_ar_payload_len   (io_outputs_2_ar_validPipe_payload_len_1[7:0]                            ), //i
    .io_inputs_1_ar_payload_size  (io_outputs_2_ar_validPipe_payload_size_1[2:0]                           ), //i
    .io_inputs_1_ar_payload_burst (io_outputs_2_ar_validPipe_payload_burst_1[1:0]                          ), //i
    .io_inputs_1_r_valid          (axi4ReadOnlyArbiter_5_io_inputs_1_r_valid                               ), //o
    .io_inputs_1_r_ready          (io_axiOut_readOnly_decoder_1_io_outputs_2_r_ready                       ), //i
    .io_inputs_1_r_payload_data   (axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_data[31:0]                  ), //o
    .io_inputs_1_r_payload_id     (axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_id[4:0]                     ), //o
    .io_inputs_1_r_payload_resp   (axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_resp[1:0]                   ), //o
    .io_inputs_1_r_payload_last   (axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_last                        ), //o
    .io_inputs_2_ar_valid         (io_outputs_2_ar_validPipe_valid_2                                       ), //i
    .io_inputs_2_ar_ready         (axi4ReadOnlyArbiter_5_io_inputs_2_ar_ready                              ), //o
    .io_inputs_2_ar_payload_addr  (io_outputs_2_ar_validPipe_payload_addr_2[31:0]                          ), //i
    .io_inputs_2_ar_payload_id    (axi4ReadOnlyArbiter_5_io_inputs_2_ar_payload_id[4:0]                    ), //i
    .io_inputs_2_ar_payload_len   (io_outputs_2_ar_validPipe_payload_len_2[7:0]                            ), //i
    .io_inputs_2_ar_payload_size  (io_outputs_2_ar_validPipe_payload_size_2[2:0]                           ), //i
    .io_inputs_2_ar_payload_burst (io_outputs_2_ar_validPipe_payload_burst_2[1:0]                          ), //i
    .io_inputs_2_r_valid          (axi4ReadOnlyArbiter_5_io_inputs_2_r_valid                               ), //o
    .io_inputs_2_r_ready          (DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_r_ready), //i
    .io_inputs_2_r_payload_data   (axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_data[31:0]                  ), //o
    .io_inputs_2_r_payload_id     (axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_id[4:0]                     ), //o
    .io_inputs_2_r_payload_resp   (axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_resp[1:0]                   ), //o
    .io_inputs_2_r_payload_last   (axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_last                        ), //o
    .io_inputs_3_ar_valid         (io_outputs_2_ar_validPipe_valid_3                                       ), //i
    .io_inputs_3_ar_ready         (axi4ReadOnlyArbiter_5_io_inputs_3_ar_ready                              ), //o
    .io_inputs_3_ar_payload_addr  (io_outputs_2_ar_validPipe_payload_addr_3[31:0]                          ), //i
    .io_inputs_3_ar_payload_id    (axi4ReadOnlyArbiter_5_io_inputs_3_ar_payload_id[4:0]                    ), //i
    .io_inputs_3_ar_payload_len   (io_outputs_2_ar_validPipe_payload_len_3[7:0]                            ), //i
    .io_inputs_3_ar_payload_size  (io_outputs_2_ar_validPipe_payload_size_3[2:0]                           ), //i
    .io_inputs_3_ar_payload_burst (io_outputs_2_ar_validPipe_payload_burst_3[1:0]                          ), //i
    .io_inputs_3_r_valid          (axi4ReadOnlyArbiter_5_io_inputs_3_r_valid                               ), //o
    .io_inputs_3_r_ready          (CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_r_ready), //i
    .io_inputs_3_r_payload_data   (axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_data[31:0]                  ), //o
    .io_inputs_3_r_payload_id     (axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_id[4:0]                     ), //o
    .io_inputs_3_r_payload_resp   (axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_resp[1:0]                   ), //o
    .io_inputs_3_r_payload_last   (axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_last                        ), //o
    .io_output_ar_valid           (axi4ReadOnlyArbiter_5_io_output_ar_valid                                ), //o
    .io_output_ar_ready           (uartAxi_ar_ready                                                        ), //i
    .io_output_ar_payload_addr    (axi4ReadOnlyArbiter_5_io_output_ar_payload_addr[31:0]                   ), //o
    .io_output_ar_payload_id      (axi4ReadOnlyArbiter_5_io_output_ar_payload_id[6:0]                      ), //o
    .io_output_ar_payload_len     (axi4ReadOnlyArbiter_5_io_output_ar_payload_len[7:0]                     ), //o
    .io_output_ar_payload_size    (axi4ReadOnlyArbiter_5_io_output_ar_payload_size[2:0]                    ), //o
    .io_output_ar_payload_burst   (axi4ReadOnlyArbiter_5_io_output_ar_payload_burst[1:0]                   ), //o
    .io_output_r_valid            (uartAxi_r_valid                                                         ), //i
    .io_output_r_ready            (axi4ReadOnlyArbiter_5_io_output_r_ready                                 ), //o
    .io_output_r_payload_data     (uartAxi_r_payload_data[31:0]                                            ), //i
    .io_output_r_payload_id       (uartAxi_r_payload_id[6:0]                                               ), //i
    .io_output_r_payload_resp     (uartAxi_r_payload_resp[1:0]                                             ), //i
    .io_output_r_payload_last     (uartAxi_r_payload_last                                                  ), //i
    .clk                          (clk                                                                     ), //i
    .reset                        (reset                                                                   )  //i
  );
  Axi4WriteOnlyArbiter axi4WriteOnlyArbiter_5 (
    .io_inputs_0_aw_valid         (io_outputs_2_aw_validPipe_valid                                                       ), //i
    .io_inputs_0_aw_ready         (axi4WriteOnlyArbiter_5_io_inputs_0_aw_ready                                           ), //o
    .io_inputs_0_aw_payload_addr  (io_outputs_2_aw_validPipe_payload_addr[31:0]                                          ), //i
    .io_inputs_0_aw_payload_id    (axi4WriteOnlyArbiter_5_io_inputs_0_aw_payload_id[4:0]                                 ), //i
    .io_inputs_0_aw_payload_len   (io_outputs_2_aw_validPipe_payload_len[7:0]                                            ), //i
    .io_inputs_0_aw_payload_size  (io_outputs_2_aw_validPipe_payload_size[2:0]                                           ), //i
    .io_inputs_0_aw_payload_burst (io_outputs_2_aw_validPipe_payload_burst[1:0]                                          ), //i
    .io_inputs_0_w_valid          (io_axiOut_writeOnly_decoder_io_outputs_2_w_valid                                      ), //i
    .io_inputs_0_w_ready          (axi4WriteOnlyArbiter_5_io_inputs_0_w_ready                                            ), //o
    .io_inputs_0_w_payload_data   (io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_data[31:0]                         ), //i
    .io_inputs_0_w_payload_strb   (io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_strb[3:0]                          ), //i
    .io_inputs_0_w_payload_last   (io_axiOut_writeOnly_decoder_io_outputs_2_w_payload_last                               ), //i
    .io_inputs_0_b_valid          (axi4WriteOnlyArbiter_5_io_inputs_0_b_valid                                            ), //o
    .io_inputs_0_b_ready          (io_axiOut_writeOnly_decoder_io_outputs_2_b_ready                                      ), //i
    .io_inputs_0_b_payload_id     (axi4WriteOnlyArbiter_5_io_inputs_0_b_payload_id[4:0]                                  ), //o
    .io_inputs_0_b_payload_resp   (axi4WriteOnlyArbiter_5_io_inputs_0_b_payload_resp[1:0]                                ), //o
    .io_inputs_1_aw_valid         (io_outputs_2_aw_validPipe_valid_1                                                     ), //i
    .io_inputs_1_aw_ready         (axi4WriteOnlyArbiter_5_io_inputs_1_aw_ready                                           ), //o
    .io_inputs_1_aw_payload_addr  (io_outputs_2_aw_validPipe_payload_addr_1[31:0]                                        ), //i
    .io_inputs_1_aw_payload_id    (axi4WriteOnlyArbiter_5_io_inputs_1_aw_payload_id[4:0]                                 ), //i
    .io_inputs_1_aw_payload_len   (io_outputs_2_aw_validPipe_payload_len_1[7:0]                                          ), //i
    .io_inputs_1_aw_payload_size  (io_outputs_2_aw_validPipe_payload_size_1[2:0]                                         ), //i
    .io_inputs_1_aw_payload_burst (io_outputs_2_aw_validPipe_payload_burst_1[1:0]                                        ), //i
    .io_inputs_1_w_valid          (io_axiOut_writeOnly_decoder_1_io_outputs_2_w_valid                                    ), //i
    .io_inputs_1_w_ready          (axi4WriteOnlyArbiter_5_io_inputs_1_w_ready                                            ), //o
    .io_inputs_1_w_payload_data   (io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_data[31:0]                       ), //i
    .io_inputs_1_w_payload_strb   (io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_strb[3:0]                        ), //i
    .io_inputs_1_w_payload_last   (io_axiOut_writeOnly_decoder_1_io_outputs_2_w_payload_last                             ), //i
    .io_inputs_1_b_valid          (axi4WriteOnlyArbiter_5_io_inputs_1_b_valid                                            ), //o
    .io_inputs_1_b_ready          (io_axiOut_writeOnly_decoder_1_io_outputs_2_b_ready                                    ), //i
    .io_inputs_1_b_payload_id     (axi4WriteOnlyArbiter_5_io_inputs_1_b_payload_id[4:0]                                  ), //o
    .io_inputs_1_b_payload_resp   (axi4WriteOnlyArbiter_5_io_inputs_1_b_payload_resp[1:0]                                ), //o
    .io_inputs_2_aw_valid         (io_outputs_2_aw_validPipe_valid_2                                                     ), //i
    .io_inputs_2_aw_ready         (axi4WriteOnlyArbiter_5_io_inputs_2_aw_ready                                           ), //o
    .io_inputs_2_aw_payload_addr  (io_outputs_2_aw_validPipe_payload_addr_2[31:0]                                        ), //i
    .io_inputs_2_aw_payload_id    (axi4WriteOnlyArbiter_5_io_inputs_2_aw_payload_id[4:0]                                 ), //i
    .io_inputs_2_aw_payload_len   (io_outputs_2_aw_validPipe_payload_len_2[7:0]                                          ), //i
    .io_inputs_2_aw_payload_size  (io_outputs_2_aw_validPipe_payload_size_2[2:0]                                         ), //i
    .io_inputs_2_aw_payload_burst (io_outputs_2_aw_validPipe_payload_burst_2[1:0]                                        ), //i
    .io_inputs_2_w_valid          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_valid             ), //i
    .io_inputs_2_w_ready          (axi4WriteOnlyArbiter_5_io_inputs_2_w_ready                                            ), //o
    .io_inputs_2_w_payload_data   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_data[31:0]), //i
    .io_inputs_2_w_payload_strb   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_strb[3:0] ), //i
    .io_inputs_2_w_payload_last   (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_w_payload_last      ), //i
    .io_inputs_2_b_valid          (axi4WriteOnlyArbiter_5_io_inputs_2_b_valid                                            ), //o
    .io_inputs_2_b_ready          (DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_b_ready             ), //i
    .io_inputs_2_b_payload_id     (axi4WriteOnlyArbiter_5_io_inputs_2_b_payload_id[4:0]                                  ), //o
    .io_inputs_2_b_payload_resp   (axi4WriteOnlyArbiter_5_io_inputs_2_b_payload_resp[1:0]                                ), //o
    .io_inputs_3_aw_valid         (io_outputs_2_aw_validPipe_valid_3                                                     ), //i
    .io_inputs_3_aw_ready         (axi4WriteOnlyArbiter_5_io_inputs_3_aw_ready                                           ), //o
    .io_inputs_3_aw_payload_addr  (io_outputs_2_aw_validPipe_payload_addr_3[31:0]                                        ), //i
    .io_inputs_3_aw_payload_id    (axi4WriteOnlyArbiter_5_io_inputs_3_aw_payload_id[4:0]                                 ), //i
    .io_inputs_3_aw_payload_len   (io_outputs_2_aw_validPipe_payload_len_3[7:0]                                          ), //i
    .io_inputs_3_aw_payload_size  (io_outputs_2_aw_validPipe_payload_size_3[2:0]                                         ), //i
    .io_inputs_3_aw_payload_burst (io_outputs_2_aw_validPipe_payload_burst_3[1:0]                                        ), //i
    .io_inputs_3_w_valid          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_valid             ), //i
    .io_inputs_3_w_ready          (axi4WriteOnlyArbiter_5_io_inputs_3_w_ready                                            ), //o
    .io_inputs_3_w_payload_data   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_data[31:0]), //i
    .io_inputs_3_w_payload_strb   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_strb[3:0] ), //i
    .io_inputs_3_w_payload_last   (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_w_payload_last      ), //i
    .io_inputs_3_b_valid          (axi4WriteOnlyArbiter_5_io_inputs_3_b_valid                                            ), //o
    .io_inputs_3_b_ready          (CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_b_ready             ), //i
    .io_inputs_3_b_payload_id     (axi4WriteOnlyArbiter_5_io_inputs_3_b_payload_id[4:0]                                  ), //o
    .io_inputs_3_b_payload_resp   (axi4WriteOnlyArbiter_5_io_inputs_3_b_payload_resp[1:0]                                ), //o
    .io_output_aw_valid           (axi4WriteOnlyArbiter_5_io_output_aw_valid                                             ), //o
    .io_output_aw_ready           (uartAxi_aw_ready                                                                      ), //i
    .io_output_aw_payload_addr    (axi4WriteOnlyArbiter_5_io_output_aw_payload_addr[31:0]                                ), //o
    .io_output_aw_payload_id      (axi4WriteOnlyArbiter_5_io_output_aw_payload_id[6:0]                                   ), //o
    .io_output_aw_payload_len     (axi4WriteOnlyArbiter_5_io_output_aw_payload_len[7:0]                                  ), //o
    .io_output_aw_payload_size    (axi4WriteOnlyArbiter_5_io_output_aw_payload_size[2:0]                                 ), //o
    .io_output_aw_payload_burst   (axi4WriteOnlyArbiter_5_io_output_aw_payload_burst[1:0]                                ), //o
    .io_output_w_valid            (axi4WriteOnlyArbiter_5_io_output_w_valid                                              ), //o
    .io_output_w_ready            (uartAxi_w_ready                                                                       ), //i
    .io_output_w_payload_data     (axi4WriteOnlyArbiter_5_io_output_w_payload_data[31:0]                                 ), //o
    .io_output_w_payload_strb     (axi4WriteOnlyArbiter_5_io_output_w_payload_strb[3:0]                                  ), //o
    .io_output_w_payload_last     (axi4WriteOnlyArbiter_5_io_output_w_payload_last                                       ), //o
    .io_output_b_valid            (uartAxi_b_valid                                                                       ), //i
    .io_output_b_ready            (axi4WriteOnlyArbiter_5_io_output_b_ready                                              ), //o
    .io_output_b_payload_id       (uartAxi_b_payload_id[6:0]                                                             ), //i
    .io_output_b_payload_resp     (uartAxi_b_payload_resp[1:0]                                                           ), //i
    .clk                          (clk                                                                                   ), //i
    .reset                        (reset                                                                                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC io_switch_btn_buffercc (
    .io_dataIn  (io_switch_btn                    ), //i
    .io_dataOut (io_switch_btn_buffercc_io_dataOut), //o
    .clk        (clk                              ), //i
    .reset      (reset                            )  //i
  );
  always @(*) begin
    case(_zz_CommitPlugin_logic_s0_committedThisCycle_comb_1)
      1'b0 : _zz_CommitPlugin_logic_s0_committedThisCycle_comb = 1'b0;
      default : _zz_CommitPlugin_logic_s0_committedThisCycle_comb = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_CommitPlugin_logic_s0_recycledThisCycle_comb_1)
      1'b0 : _zz_CommitPlugin_logic_s0_recycledThisCycle_comb = 1'b0;
      default : _zz_CommitPlugin_logic_s0_recycledThisCycle_comb = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_DispatchPlugin_logic_destinationIqReady_4)
      2'b00 : _zz_DispatchPlugin_logic_destinationIqReady_3 = DispatchPlugin_logic_iqRegs_0_1_ready;
      2'b01 : _zz_DispatchPlugin_logic_destinationIqReady_3 = DispatchPlugin_logic_iqRegs_1_1_ready;
      2'b10 : _zz_DispatchPlugin_logic_destinationIqReady_3 = DispatchPlugin_logic_iqRegs_2_1_ready;
      default : _zz_DispatchPlugin_logic_destinationIqReady_3 = DispatchPlugin_logic_iqRegs_3_1_ready;
    endcase
  end

  always @(*) begin
    case(AluIntEU_AluIntEuPlugin_gprReadPorts_0_address)
      6'b000000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_0;
      6'b000001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_1;
      6'b000010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_2;
      6'b000011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_3;
      6'b000100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_4;
      6'b000101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_5;
      6'b000110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_6;
      6'b000111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_7;
      6'b001000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_8;
      6'b001001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_9;
      6'b001010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_10;
      6'b001011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_11;
      6'b001100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_12;
      6'b001101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_13;
      6'b001110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_14;
      6'b001111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_15;
      6'b010000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_16;
      6'b010001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_17;
      6'b010010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_18;
      6'b010011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_19;
      6'b010100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_20;
      6'b010101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_21;
      6'b010110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_22;
      6'b010111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_23;
      6'b011000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_24;
      6'b011001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_25;
      6'b011010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_26;
      6'b011011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_27;
      6'b011100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_28;
      6'b011101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_29;
      6'b011110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_30;
      6'b011111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_31;
      6'b100000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_32;
      6'b100001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_33;
      6'b100010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_34;
      6'b100011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_35;
      6'b100100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_36;
      6'b100101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_37;
      6'b100110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_38;
      6'b100111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_39;
      6'b101000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_40;
      6'b101001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_41;
      6'b101010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_42;
      6'b101011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_43;
      6'b101100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_44;
      6'b101101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_45;
      6'b101110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_46;
      6'b101111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_47;
      6'b110000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_48;
      6'b110001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_49;
      6'b110010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_50;
      6'b110011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_51;
      6'b110100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_52;
      6'b110101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_53;
      6'b110110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_54;
      6'b110111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_55;
      6'b111000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_56;
      6'b111001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_57;
      6'b111010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_58;
      6'b111011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_59;
      6'b111100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_60;
      6'b111101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_61;
      6'b111110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_62;
      default : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_63;
    endcase
  end

  always @(*) begin
    case(AluIntEU_AluIntEuPlugin_gprReadPorts_1_address)
      6'b000000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_0;
      6'b000001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_1;
      6'b000010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_2;
      6'b000011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_3;
      6'b000100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_4;
      6'b000101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_5;
      6'b000110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_6;
      6'b000111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_7;
      6'b001000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_8;
      6'b001001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_9;
      6'b001010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_10;
      6'b001011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_11;
      6'b001100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_12;
      6'b001101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_13;
      6'b001110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_14;
      6'b001111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_15;
      6'b010000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_16;
      6'b010001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_17;
      6'b010010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_18;
      6'b010011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_19;
      6'b010100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_20;
      6'b010101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_21;
      6'b010110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_22;
      6'b010111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_23;
      6'b011000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_24;
      6'b011001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_25;
      6'b011010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_26;
      6'b011011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_27;
      6'b011100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_28;
      6'b011101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_29;
      6'b011110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_30;
      6'b011111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_31;
      6'b100000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_32;
      6'b100001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_33;
      6'b100010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_34;
      6'b100011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_35;
      6'b100100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_36;
      6'b100101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_37;
      6'b100110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_38;
      6'b100111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_39;
      6'b101000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_40;
      6'b101001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_41;
      6'b101010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_42;
      6'b101011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_43;
      6'b101100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_44;
      6'b101101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_45;
      6'b101110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_46;
      6'b101111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_47;
      6'b110000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_48;
      6'b110001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_49;
      6'b110010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_50;
      6'b110011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_51;
      6'b110100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_52;
      6'b110101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_53;
      6'b110110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_54;
      6'b110111 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_55;
      6'b111000 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_56;
      6'b111001 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_57;
      6'b111010 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_58;
      6'b111011 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_59;
      6'b111100 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_60;
      6'b111101 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_61;
      6'b111110 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_62;
      default : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_63;
    endcase
  end

  always @(*) begin
    case(MulEU_MulEuPlugin_gprReadPorts_0_address)
      6'b000000 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_0;
      6'b000001 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_1;
      6'b000010 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_2;
      6'b000011 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_3;
      6'b000100 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_4;
      6'b000101 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_5;
      6'b000110 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_6;
      6'b000111 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_7;
      6'b001000 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_8;
      6'b001001 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_9;
      6'b001010 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_10;
      6'b001011 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_11;
      6'b001100 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_12;
      6'b001101 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_13;
      6'b001110 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_14;
      6'b001111 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_15;
      6'b010000 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_16;
      6'b010001 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_17;
      6'b010010 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_18;
      6'b010011 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_19;
      6'b010100 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_20;
      6'b010101 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_21;
      6'b010110 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_22;
      6'b010111 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_23;
      6'b011000 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_24;
      6'b011001 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_25;
      6'b011010 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_26;
      6'b011011 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_27;
      6'b011100 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_28;
      6'b011101 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_29;
      6'b011110 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_30;
      6'b011111 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_31;
      6'b100000 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_32;
      6'b100001 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_33;
      6'b100010 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_34;
      6'b100011 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_35;
      6'b100100 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_36;
      6'b100101 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_37;
      6'b100110 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_38;
      6'b100111 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_39;
      6'b101000 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_40;
      6'b101001 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_41;
      6'b101010 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_42;
      6'b101011 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_43;
      6'b101100 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_44;
      6'b101101 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_45;
      6'b101110 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_46;
      6'b101111 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_47;
      6'b110000 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_48;
      6'b110001 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_49;
      6'b110010 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_50;
      6'b110011 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_51;
      6'b110100 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_52;
      6'b110101 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_53;
      6'b110110 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_54;
      6'b110111 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_55;
      6'b111000 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_56;
      6'b111001 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_57;
      6'b111010 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_58;
      6'b111011 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_59;
      6'b111100 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_60;
      6'b111101 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_61;
      6'b111110 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_62;
      default : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_63;
    endcase
  end

  always @(*) begin
    case(MulEU_MulEuPlugin_gprReadPorts_1_address)
      6'b000000 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_0;
      6'b000001 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_1;
      6'b000010 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_2;
      6'b000011 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_3;
      6'b000100 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_4;
      6'b000101 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_5;
      6'b000110 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_6;
      6'b000111 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_7;
      6'b001000 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_8;
      6'b001001 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_9;
      6'b001010 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_10;
      6'b001011 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_11;
      6'b001100 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_12;
      6'b001101 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_13;
      6'b001110 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_14;
      6'b001111 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_15;
      6'b010000 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_16;
      6'b010001 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_17;
      6'b010010 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_18;
      6'b010011 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_19;
      6'b010100 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_20;
      6'b010101 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_21;
      6'b010110 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_22;
      6'b010111 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_23;
      6'b011000 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_24;
      6'b011001 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_25;
      6'b011010 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_26;
      6'b011011 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_27;
      6'b011100 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_28;
      6'b011101 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_29;
      6'b011110 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_30;
      6'b011111 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_31;
      6'b100000 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_32;
      6'b100001 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_33;
      6'b100010 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_34;
      6'b100011 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_35;
      6'b100100 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_36;
      6'b100101 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_37;
      6'b100110 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_38;
      6'b100111 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_39;
      6'b101000 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_40;
      6'b101001 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_41;
      6'b101010 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_42;
      6'b101011 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_43;
      6'b101100 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_44;
      6'b101101 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_45;
      6'b101110 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_46;
      6'b101111 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_47;
      6'b110000 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_48;
      6'b110001 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_49;
      6'b110010 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_50;
      6'b110011 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_51;
      6'b110100 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_52;
      6'b110101 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_53;
      6'b110110 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_54;
      6'b110111 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_55;
      6'b111000 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_56;
      6'b111001 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_57;
      6'b111010 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_58;
      6'b111011 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_59;
      6'b111100 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_60;
      6'b111101 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_61;
      6'b111110 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_62;
      default : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_63;
    endcase
  end

  always @(*) begin
    case(BranchEU_BranchEuPlugin_gprReadPorts_0_address)
      6'b000000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_0;
      6'b000001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_1;
      6'b000010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_2;
      6'b000011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_3;
      6'b000100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_4;
      6'b000101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_5;
      6'b000110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_6;
      6'b000111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_7;
      6'b001000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_8;
      6'b001001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_9;
      6'b001010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_10;
      6'b001011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_11;
      6'b001100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_12;
      6'b001101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_13;
      6'b001110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_14;
      6'b001111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_15;
      6'b010000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_16;
      6'b010001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_17;
      6'b010010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_18;
      6'b010011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_19;
      6'b010100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_20;
      6'b010101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_21;
      6'b010110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_22;
      6'b010111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_23;
      6'b011000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_24;
      6'b011001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_25;
      6'b011010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_26;
      6'b011011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_27;
      6'b011100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_28;
      6'b011101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_29;
      6'b011110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_30;
      6'b011111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_31;
      6'b100000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_32;
      6'b100001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_33;
      6'b100010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_34;
      6'b100011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_35;
      6'b100100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_36;
      6'b100101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_37;
      6'b100110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_38;
      6'b100111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_39;
      6'b101000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_40;
      6'b101001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_41;
      6'b101010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_42;
      6'b101011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_43;
      6'b101100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_44;
      6'b101101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_45;
      6'b101110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_46;
      6'b101111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_47;
      6'b110000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_48;
      6'b110001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_49;
      6'b110010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_50;
      6'b110011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_51;
      6'b110100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_52;
      6'b110101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_53;
      6'b110110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_54;
      6'b110111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_55;
      6'b111000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_56;
      6'b111001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_57;
      6'b111010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_58;
      6'b111011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_59;
      6'b111100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_60;
      6'b111101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_61;
      6'b111110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_62;
      default : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = PhysicalRegFilePlugin_logic_regFile_63;
    endcase
  end

  always @(*) begin
    case(BranchEU_BranchEuPlugin_gprReadPorts_1_address)
      6'b000000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_0;
      6'b000001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_1;
      6'b000010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_2;
      6'b000011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_3;
      6'b000100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_4;
      6'b000101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_5;
      6'b000110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_6;
      6'b000111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_7;
      6'b001000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_8;
      6'b001001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_9;
      6'b001010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_10;
      6'b001011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_11;
      6'b001100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_12;
      6'b001101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_13;
      6'b001110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_14;
      6'b001111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_15;
      6'b010000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_16;
      6'b010001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_17;
      6'b010010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_18;
      6'b010011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_19;
      6'b010100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_20;
      6'b010101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_21;
      6'b010110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_22;
      6'b010111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_23;
      6'b011000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_24;
      6'b011001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_25;
      6'b011010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_26;
      6'b011011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_27;
      6'b011100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_28;
      6'b011101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_29;
      6'b011110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_30;
      6'b011111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_31;
      6'b100000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_32;
      6'b100001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_33;
      6'b100010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_34;
      6'b100011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_35;
      6'b100100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_36;
      6'b100101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_37;
      6'b100110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_38;
      6'b100111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_39;
      6'b101000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_40;
      6'b101001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_41;
      6'b101010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_42;
      6'b101011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_43;
      6'b101100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_44;
      6'b101101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_45;
      6'b101110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_46;
      6'b101111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_47;
      6'b110000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_48;
      6'b110001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_49;
      6'b110010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_50;
      6'b110011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_51;
      6'b110100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_52;
      6'b110101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_53;
      6'b110110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_54;
      6'b110111 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_55;
      6'b111000 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_56;
      6'b111001 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_57;
      6'b111010 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_58;
      6'b111011 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_59;
      6'b111100 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_60;
      6'b111101 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_61;
      6'b111110 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_62;
      default : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = PhysicalRegFilePlugin_logic_regFile_63;
    endcase
  end

  always @(*) begin
    case(LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_address)
      6'b000000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_0;
      6'b000001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_1;
      6'b000010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_2;
      6'b000011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_3;
      6'b000100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_4;
      6'b000101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_5;
      6'b000110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_6;
      6'b000111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_7;
      6'b001000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_8;
      6'b001001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_9;
      6'b001010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_10;
      6'b001011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_11;
      6'b001100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_12;
      6'b001101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_13;
      6'b001110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_14;
      6'b001111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_15;
      6'b010000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_16;
      6'b010001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_17;
      6'b010010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_18;
      6'b010011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_19;
      6'b010100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_20;
      6'b010101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_21;
      6'b010110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_22;
      6'b010111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_23;
      6'b011000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_24;
      6'b011001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_25;
      6'b011010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_26;
      6'b011011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_27;
      6'b011100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_28;
      6'b011101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_29;
      6'b011110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_30;
      6'b011111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_31;
      6'b100000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_32;
      6'b100001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_33;
      6'b100010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_34;
      6'b100011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_35;
      6'b100100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_36;
      6'b100101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_37;
      6'b100110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_38;
      6'b100111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_39;
      6'b101000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_40;
      6'b101001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_41;
      6'b101010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_42;
      6'b101011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_43;
      6'b101100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_44;
      6'b101101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_45;
      6'b101110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_46;
      6'b101111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_47;
      6'b110000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_48;
      6'b110001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_49;
      6'b110010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_50;
      6'b110011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_51;
      6'b110100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_52;
      6'b110101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_53;
      6'b110110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_54;
      6'b110111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_55;
      6'b111000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_56;
      6'b111001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_57;
      6'b111010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_58;
      6'b111011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_59;
      6'b111100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_60;
      6'b111101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_61;
      6'b111110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_62;
      default : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = PhysicalRegFilePlugin_logic_regFile_63;
    endcase
  end

  always @(*) begin
    case(LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_address)
      6'b000000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_0;
      6'b000001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_1;
      6'b000010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_2;
      6'b000011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_3;
      6'b000100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_4;
      6'b000101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_5;
      6'b000110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_6;
      6'b000111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_7;
      6'b001000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_8;
      6'b001001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_9;
      6'b001010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_10;
      6'b001011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_11;
      6'b001100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_12;
      6'b001101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_13;
      6'b001110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_14;
      6'b001111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_15;
      6'b010000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_16;
      6'b010001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_17;
      6'b010010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_18;
      6'b010011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_19;
      6'b010100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_20;
      6'b010101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_21;
      6'b010110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_22;
      6'b010111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_23;
      6'b011000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_24;
      6'b011001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_25;
      6'b011010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_26;
      6'b011011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_27;
      6'b011100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_28;
      6'b011101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_29;
      6'b011110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_30;
      6'b011111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_31;
      6'b100000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_32;
      6'b100001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_33;
      6'b100010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_34;
      6'b100011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_35;
      6'b100100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_36;
      6'b100101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_37;
      6'b100110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_38;
      6'b100111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_39;
      6'b101000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_40;
      6'b101001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_41;
      6'b101010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_42;
      6'b101011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_43;
      6'b101100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_44;
      6'b101101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_45;
      6'b101110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_46;
      6'b101111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_47;
      6'b110000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_48;
      6'b110001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_49;
      6'b110010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_50;
      6'b110011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_51;
      6'b110100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_52;
      6'b110101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_53;
      6'b110110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_54;
      6'b110111 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_55;
      6'b111000 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_56;
      6'b111001 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_57;
      6'b111010 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_58;
      6'b111011 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_59;
      6'b111100 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_60;
      6'b111101 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_61;
      6'b111110 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_62;
      default : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = PhysicalRegFilePlugin_logic_regFile_63;
    endcase
  end

  always @(*) begin
    case(FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_startInstructionIndex)
      2'b00 : _zz__zz_71 = FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_0_isBranch;
      2'b01 : _zz__zz_71 = FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_1_isBranch;
      2'b10 : _zz__zz_71 = FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_2_isBranch;
      default : _zz__zz_71 = FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_predecodeInfos_3_isBranch;
    endcase
  end

  always @(*) begin
    case(ICachePlugin_logic_pipeline_f1_f1_index)
      7'b0000000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_0_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_0_1;
      end
      7'b0000001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_1_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_1_1;
      end
      7'b0000010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_2_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_2_1;
      end
      7'b0000011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_3_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_3_1;
      end
      7'b0000100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_4_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_4_1;
      end
      7'b0000101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_5_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_5_1;
      end
      7'b0000110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_6_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_6_1;
      end
      7'b0000111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_7_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_7_1;
      end
      7'b0001000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_8_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_8_1;
      end
      7'b0001001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_9_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_9_1;
      end
      7'b0001010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_10_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_10_1;
      end
      7'b0001011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_11_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_11_1;
      end
      7'b0001100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_12_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_12_1;
      end
      7'b0001101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_13_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_13_1;
      end
      7'b0001110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_14_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_14_1;
      end
      7'b0001111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_15_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_15_1;
      end
      7'b0010000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_16_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_16_1;
      end
      7'b0010001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_17_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_17_1;
      end
      7'b0010010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_18_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_18_1;
      end
      7'b0010011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_19_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_19_1;
      end
      7'b0010100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_20_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_20_1;
      end
      7'b0010101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_21_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_21_1;
      end
      7'b0010110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_22_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_22_1;
      end
      7'b0010111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_23_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_23_1;
      end
      7'b0011000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_24_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_24_1;
      end
      7'b0011001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_25_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_25_1;
      end
      7'b0011010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_26_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_26_1;
      end
      7'b0011011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_27_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_27_1;
      end
      7'b0011100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_28_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_28_1;
      end
      7'b0011101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_29_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_29_1;
      end
      7'b0011110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_30_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_30_1;
      end
      7'b0011111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_31_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_31_1;
      end
      7'b0100000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_32_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_32_1;
      end
      7'b0100001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_33_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_33_1;
      end
      7'b0100010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_34_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_34_1;
      end
      7'b0100011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_35_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_35_1;
      end
      7'b0100100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_36_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_36_1;
      end
      7'b0100101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_37_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_37_1;
      end
      7'b0100110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_38_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_38_1;
      end
      7'b0100111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_39_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_39_1;
      end
      7'b0101000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_40_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_40_1;
      end
      7'b0101001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_41_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_41_1;
      end
      7'b0101010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_42_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_42_1;
      end
      7'b0101011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_43_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_43_1;
      end
      7'b0101100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_44_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_44_1;
      end
      7'b0101101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_45_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_45_1;
      end
      7'b0101110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_46_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_46_1;
      end
      7'b0101111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_47_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_47_1;
      end
      7'b0110000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_48_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_48_1;
      end
      7'b0110001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_49_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_49_1;
      end
      7'b0110010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_50_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_50_1;
      end
      7'b0110011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_51_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_51_1;
      end
      7'b0110100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_52_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_52_1;
      end
      7'b0110101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_53_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_53_1;
      end
      7'b0110110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_54_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_54_1;
      end
      7'b0110111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_55_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_55_1;
      end
      7'b0111000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_56_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_56_1;
      end
      7'b0111001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_57_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_57_1;
      end
      7'b0111010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_58_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_58_1;
      end
      7'b0111011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_59_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_59_1;
      end
      7'b0111100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_60_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_60_1;
      end
      7'b0111101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_61_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_61_1;
      end
      7'b0111110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_62_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_62_1;
      end
      7'b0111111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_63_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_63_1;
      end
      7'b1000000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_64_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_64_1;
      end
      7'b1000001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_65_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_65_1;
      end
      7'b1000010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_66_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_66_1;
      end
      7'b1000011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_67_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_67_1;
      end
      7'b1000100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_68_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_68_1;
      end
      7'b1000101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_69_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_69_1;
      end
      7'b1000110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_70_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_70_1;
      end
      7'b1000111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_71_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_71_1;
      end
      7'b1001000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_72_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_72_1;
      end
      7'b1001001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_73_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_73_1;
      end
      7'b1001010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_74_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_74_1;
      end
      7'b1001011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_75_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_75_1;
      end
      7'b1001100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_76_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_76_1;
      end
      7'b1001101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_77_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_77_1;
      end
      7'b1001110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_78_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_78_1;
      end
      7'b1001111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_79_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_79_1;
      end
      7'b1010000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_80_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_80_1;
      end
      7'b1010001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_81_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_81_1;
      end
      7'b1010010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_82_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_82_1;
      end
      7'b1010011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_83_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_83_1;
      end
      7'b1010100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_84_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_84_1;
      end
      7'b1010101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_85_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_85_1;
      end
      7'b1010110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_86_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_86_1;
      end
      7'b1010111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_87_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_87_1;
      end
      7'b1011000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_88_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_88_1;
      end
      7'b1011001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_89_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_89_1;
      end
      7'b1011010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_90_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_90_1;
      end
      7'b1011011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_91_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_91_1;
      end
      7'b1011100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_92_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_92_1;
      end
      7'b1011101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_93_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_93_1;
      end
      7'b1011110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_94_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_94_1;
      end
      7'b1011111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_95_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_95_1;
      end
      7'b1100000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_96_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_96_1;
      end
      7'b1100001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_97_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_97_1;
      end
      7'b1100010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_98_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_98_1;
      end
      7'b1100011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_99_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_99_1;
      end
      7'b1100100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_100_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_100_1;
      end
      7'b1100101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_101_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_101_1;
      end
      7'b1100110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_102_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_102_1;
      end
      7'b1100111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_103_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_103_1;
      end
      7'b1101000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_104_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_104_1;
      end
      7'b1101001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_105_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_105_1;
      end
      7'b1101010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_106_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_106_1;
      end
      7'b1101011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_107_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_107_1;
      end
      7'b1101100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_108_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_108_1;
      end
      7'b1101101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_109_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_109_1;
      end
      7'b1101110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_110_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_110_1;
      end
      7'b1101111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_111_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_111_1;
      end
      7'b1110000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_112_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_112_1;
      end
      7'b1110001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_113_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_113_1;
      end
      7'b1110010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_114_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_114_1;
      end
      7'b1110011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_115_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_115_1;
      end
      7'b1110100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_116_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_116_1;
      end
      7'b1110101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_117_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_117_1;
      end
      7'b1110110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_118_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_118_1;
      end
      7'b1110111 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_119_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_119_1;
      end
      7'b1111000 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_120_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_120_1;
      end
      7'b1111001 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_121_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_121_1;
      end
      7'b1111010 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_122_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_122_1;
      end
      7'b1111011 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_123_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_123_1;
      end
      7'b1111100 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_124_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_124_1;
      end
      7'b1111101 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_125_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_125_1;
      end
      7'b1111110 : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_126_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_126_1;
      end
      default : begin
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = ICachePlugin_logic_storage_valids_127_0;
        _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = ICachePlugin_logic_storage_valids_127_1;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition)
      BranchCondition_NUL : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LA_CF_FALSE";
      default : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1)
      BranchCondition_NUL : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "NUL        ";
      BranchCondition_EQ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "EQ         ";
      BranchCondition_NE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "NE         ";
      BranchCondition_LT : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "LT         ";
      BranchCondition_GE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "GE         ";
      BranchCondition_LTU : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "LTU        ";
      BranchCondition_GEU : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "GEU        ";
      BranchCondition_EQZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "EQZ        ";
      BranchCondition_NEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "NEZ        ";
      BranchCondition_LTZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "LTZ        ";
      BranchCondition_GEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "GEZ        ";
      BranchCondition_GTZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "GTZ        ";
      BranchCondition_LEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "F_NE       ";
      BranchCondition_F_LT : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "F_LT       ";
      BranchCondition_F_LE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "F_LE       ";
      BranchCondition_F_UN : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "LA_CF_FALSE";
      default : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1)
      ArchRegType_GPR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1_string = "GPR  ";
      ArchRegType_FPR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1_string = "FPR  ";
      ArchRegType_CSR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1_string = "CSR  ";
      ArchRegType_LA_CF : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1_string = "LA_CF";
      default : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2)
      BranchCondition_NUL : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "NUL        ";
      BranchCondition_EQ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "EQ         ";
      BranchCondition_NE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "NE         ";
      BranchCondition_LT : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "LT         ";
      BranchCondition_GE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "GE         ";
      BranchCondition_LTU : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "LTU        ";
      BranchCondition_GEU : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "GEU        ";
      BranchCondition_EQZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "EQZ        ";
      BranchCondition_NEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "NEZ        ";
      BranchCondition_LTZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "LTZ        ";
      BranchCondition_GEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "GEZ        ";
      BranchCondition_GTZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "GTZ        ";
      BranchCondition_LEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "F_NE       ";
      BranchCondition_F_LT : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "F_LT       ";
      BranchCondition_F_LE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "F_LE       ";
      BranchCondition_F_UN : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "LA_CF_FALSE";
      default : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2)
      ArchRegType_GPR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2_string = "GPR  ";
      ArchRegType_FPR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2_string = "FPR  ";
      ArchRegType_CSR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2_string = "CSR  ";
      ArchRegType_LA_CF : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2_string = "LA_CF";
      default : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3)
      BranchCondition_NUL : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "NUL        ";
      BranchCondition_EQ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "EQ         ";
      BranchCondition_NE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "NE         ";
      BranchCondition_LT : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "LT         ";
      BranchCondition_GE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "GE         ";
      BranchCondition_LTU : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "LTU        ";
      BranchCondition_GEU : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "GEU        ";
      BranchCondition_EQZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "EQZ        ";
      BranchCondition_NEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "NEZ        ";
      BranchCondition_LTZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "LTZ        ";
      BranchCondition_GEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "GEZ        ";
      BranchCondition_GTZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "GTZ        ";
      BranchCondition_LEZ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "F_NE       ";
      BranchCondition_F_LT : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "F_LT       ";
      BranchCondition_F_LE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "F_LE       ";
      BranchCondition_F_UN : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "LA_CF_FALSE";
      default : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3)
      ArchRegType_GPR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3_string = "GPR  ";
      ArchRegType_FPR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3_string = "FPR  ";
      ArchRegType_CSR : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3_string = "CSR  ";
      ArchRegType_LA_CF : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3_string = "LA_CF";
      default : _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode)
      IntAluExceptionCode_NONE : _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_string = "NONE            ";
      IntAluExceptionCode_UNDEFINED_ALU_OP : _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_string = "UNDEFINED_ALU_OP";
      default : _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp)
      LogicOp_NONE : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "XOR_1";
      default : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage)
      ImmUsageType_NONE : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "JUMP_OFFSET  ";
      default : _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_1)
      IntAluExceptionCode_NONE : _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_1_string = "NONE            ";
      IntAluExceptionCode_UNDEFINED_ALU_OP : _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_1_string = "UNDEFINED_ALU_OP";
      default : _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_1_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_iqEntryIn_payload_aluCtrl_logicOp)
      LogicOp_NONE : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_string = "XOR_1";
      default : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_iqEntryIn_payload_immUsage)
      ImmUsageType_NONE : _zz_io_iqEntryIn_payload_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_io_iqEntryIn_payload_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_io_iqEntryIn_payload_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_io_iqEntryIn_payload_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_io_iqEntryIn_payload_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_io_iqEntryIn_payload_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_io_iqEntryIn_payload_immUsage_string = "JUMP_OFFSET  ";
      default : _zz_io_iqEntryIn_payload_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_iqEntryIn_payload_aluCtrl_logicOp_1)
      LogicOp_NONE : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1_string = "NONE ";
      LogicOp_AND_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1_string = "AND_1";
      LogicOp_OR_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1_string = "XOR_1";
      default : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_iqEntryIn_payload_immUsage_1)
      ImmUsageType_NONE : _zz_io_iqEntryIn_payload_immUsage_1_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_io_iqEntryIn_payload_immUsage_1_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_io_iqEntryIn_payload_immUsage_1_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_io_iqEntryIn_payload_immUsage_1_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_io_iqEntryIn_payload_immUsage_1_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_io_iqEntryIn_payload_immUsage_1_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_io_iqEntryIn_payload_immUsage_1_string = "JUMP_OFFSET  ";
      default : _zz_io_iqEntryIn_payload_immUsage_1_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_iqEntryIn_payload_aluCtrl_logicOp_2)
      LogicOp_NONE : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2_string = "NONE ";
      LogicOp_AND_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2_string = "AND_1";
      LogicOp_OR_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2_string = "XOR_1";
      default : _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_iqEntryIn_payload_immUsage_2)
      ImmUsageType_NONE : _zz_io_iqEntryIn_payload_immUsage_2_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_io_iqEntryIn_payload_immUsage_2_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_io_iqEntryIn_payload_immUsage_2_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_io_iqEntryIn_payload_immUsage_2_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_io_iqEntryIn_payload_immUsage_2_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_io_iqEntryIn_payload_immUsage_2_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_io_iqEntryIn_payload_immUsage_2_string = "JUMP_OFFSET  ";
      default : _zz_io_iqEntryIn_payload_immUsage_2_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode)
      BaseUopCode_NOP : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "IDLE       ";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit)
      ExeUnitType_NONE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa)
      IsaType_UNKNOWN : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "LOONGARCH";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage)
      ImmUsageType_NONE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp)
      LogicOp_NONE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition)
      BranchCondition_NUL : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "OK          ";
      default : s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode)
      BaseUopCode_NOP : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "IDLE       ";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit)
      ExeUnitType_NONE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa)
      IsaType_UNKNOWN : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa_string = "LOONGARCH";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage)
      ImmUsageType_NONE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp)
      LogicOp_NONE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition)
      BranchCondition_NUL : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode_string = "OK          ";
      default : s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode)
      BaseUopCode_NOP : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "MUL        ";
      BaseUopCode_DIV : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "IDLE       ";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit)
      ExeUnitType_NONE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "FPU_DIV_SQRT       ";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa)
      IsaType_UNKNOWN : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "UNKNOWN  ";
      IsaType_DEMO : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "DEMO     ";
      IsaType_RISCV : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "RISCV    ";
      IsaType_LOONGARCH : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "LOONGARCH";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage)
      ImmUsageType_NONE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "JUMP_OFFSET  ";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp)
      LogicOp_NONE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "XOR_1";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition)
      BranchCondition_NUL : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LA_CF_FALSE";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest)
      MemAccessSize_B : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "D";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode)
      DecodeExCode_INVALID : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "OK          ";
      default : s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode)
      BaseUopCode_NOP : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "MUL        ";
      BaseUopCode_DIV : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "IDLE       ";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit)
      ExeUnitType_NONE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "FPU_DIV_SQRT       ";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa)
      IsaType_UNKNOWN : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "UNKNOWN  ";
      IsaType_DEMO : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "DEMO     ";
      IsaType_RISCV : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "RISCV    ";
      IsaType_LOONGARCH : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "LOONGARCH";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype)
      ArchRegType_GPR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "LA_CF";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype)
      ArchRegType_GPR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "LA_CF";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype)
      ArchRegType_GPR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "LA_CF";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage)
      ImmUsageType_NONE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "JUMP_OFFSET  ";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp)
      LogicOp_NONE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "XOR_1";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size)
      MemAccessSize_B : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "B";
      MemAccessSize_H : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "H";
      MemAccessSize_W : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "W";
      MemAccessSize_D : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "D";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition)
      BranchCondition_NUL : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LA_CF_FALSE";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "D";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "D";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest)
      MemAccessSize_B : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "D";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode)
      DecodeExCode_INVALID : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "OK          ";
      default : s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode)
      BaseUopCode_NOP : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "IDLE       ";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit)
      ExeUnitType_NONE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa)
      IsaType_UNKNOWN : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "LOONGARCH";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype)
      ArchRegType_GPR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "LA_CF";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype)
      ArchRegType_GPR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "LA_CF";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype)
      ArchRegType_GPR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "LA_CF";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage)
      ImmUsageType_NONE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp)
      LogicOp_NONE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size)
      MemAccessSize_B : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "D";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition)
      BranchCondition_NUL : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "OK          ";
      default : s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode)
      BaseUopCode_NOP : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "MUL        ";
      BaseUopCode_DIV : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "IDLE       ";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit)
      ExeUnitType_NONE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "FPU_DIV_SQRT       ";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa)
      IsaType_UNKNOWN : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "UNKNOWN  ";
      IsaType_DEMO : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "DEMO     ";
      IsaType_RISCV : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "RISCV    ";
      IsaType_LOONGARCH : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "LOONGARCH";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype)
      ArchRegType_GPR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "LA_CF";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype)
      ArchRegType_GPR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "LA_CF";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype)
      ArchRegType_GPR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "LA_CF";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage)
      ImmUsageType_NONE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "JUMP_OFFSET  ";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp)
      LogicOp_NONE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "XOR_1";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size)
      MemAccessSize_B : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "B";
      MemAccessSize_H : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "H";
      MemAccessSize_W : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "W";
      MemAccessSize_D : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "D";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition)
      BranchCondition_NUL : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "LA_CF_FALSE";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "D";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "D";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest)
      MemAccessSize_B : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "D";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode)
      DecodeExCode_INVALID : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "OK          ";
      default : s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(ROBPlugin_aggregatedFlushSignal_payload_reason)
      FlushReason_NONE : ROBPlugin_aggregatedFlushSignal_payload_reason_string = "NONE               ";
      FlushReason_FULL_FLUSH : ROBPlugin_aggregatedFlushSignal_payload_reason_string = "FULL_FLUSH         ";
      FlushReason_ROLLBACK_TO_ROB_IDX : ROBPlugin_aggregatedFlushSignal_payload_reason_string = "ROLLBACK_TO_ROB_IDX";
      default : ROBPlugin_aggregatedFlushSignal_payload_reason_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp)
      LogicOp_NONE : AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "XOR_1";
      default : AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(AluIntEU_AluIntEuPlugin_euResult_uop_immUsage)
      ImmUsageType_NONE : AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "JUMP_OFFSET  ";
      default : AluIntEU_AluIntEuPlugin_euResult_uop_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_0_0)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_0_0_0_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_0_0_0_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_0_0_0_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_0_0_0_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_0_0_0_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_0_0_0_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_0_0_0_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_0_0_0_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_0_0_0_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_0_0_0_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_0_0_0_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_0_0_0_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_0_0_0_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_0_0_0_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_0_0_0_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_0_0_0_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_0_0_0_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_0_0_0_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_0_0_0_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_0_0_0_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_0_0_0_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_0_0_0_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_0_0_0_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_0_0_0_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_0_0_0_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_0_1)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_0_0_1_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_0_0_1_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_0_0_1_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_0_0_1_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_0_0_1_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_0_0_1_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_0_0_1_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_0_0_1_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_0_0_1_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_0_0_1_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_0_0_1_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_0_0_1_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_0_0_1_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_0_0_1_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_0_0_1_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_0_0_1_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_0_0_1_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_0_0_1_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_0_0_1_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_0_0_1_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_0_0_1_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_0_0_1_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_0_0_1_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_0_0_1_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_0_0_1_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_0_2)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_0_0_2_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_0_0_2_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_0_0_2_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_0_0_2_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_0_0_2_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_0_0_2_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_0_0_2_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_0_0_2_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_0_0_2_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_0_0_2_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_0_0_2_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_0_0_2_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_0_0_2_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_0_0_2_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_0_0_2_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_0_0_2_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_0_0_2_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_0_0_2_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_0_0_2_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_0_0_2_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_0_0_2_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_0_0_2_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_0_0_2_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_0_0_2_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_0_0_2_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_0_3)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_0_0_3_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_0_0_3_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_0_0_3_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_0_0_3_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_0_0_3_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_0_0_3_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_0_0_3_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_0_0_3_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_0_0_3_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_0_0_3_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_0_0_3_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_0_0_3_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_0_0_3_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_0_0_3_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_0_0_3_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_0_0_3_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_0_0_3_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_0_0_3_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_0_0_3_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_0_0_3_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_0_0_3_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_0_0_3_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_0_0_3_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_0_0_3_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_0_0_3_string = "???????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode)
      BaseUopCode_NOP : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "IDLE       ";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit)
      ExeUnitType_NONE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa)
      IsaType_UNKNOWN : MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa_string = "LOONGARCH";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype)
      ArchRegType_GPR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype_string = "LA_CF";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage)
      ImmUsageType_NONE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size)
      MemAccessSize_B : MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size_string = "D";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_0_0)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_1_0_0_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_1_0_0_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_1_0_0_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_1_0_0_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_1_0_0_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_1_0_0_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_1_0_0_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_1_0_0_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_1_0_0_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_1_0_0_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_1_0_0_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_1_0_0_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_1_0_0_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_1_0_0_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_1_0_0_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_1_0_0_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_1_0_0_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_1_0_0_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_1_0_0_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_1_0_0_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_1_0_0_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_1_0_0_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_1_0_0_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_1_0_0_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_1_0_0_string = "???????????";
    endcase
  end
  always @(*) begin
    case(BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition)
      BranchCondition_NUL : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "LA_CF_FALSE";
      default : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_0_0)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_2_0_0_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_2_0_0_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_2_0_0_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_2_0_0_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_2_0_0_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_2_0_0_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_2_0_0_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_2_0_0_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_2_0_0_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_2_0_0_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_2_0_0_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_2_0_0_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_2_0_0_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_2_0_0_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_2_0_0_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_2_0_0_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_2_0_0_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_2_0_0_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_2_0_0_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_2_0_0_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_2_0_0_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_2_0_0_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_2_0_0_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_2_0_0_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_2_0_0_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_0_1)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_2_0_1_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_2_0_1_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_2_0_1_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_2_0_1_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_2_0_1_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_2_0_1_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_2_0_1_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_2_0_1_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_2_0_1_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_2_0_1_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_2_0_1_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_2_0_1_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_2_0_1_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_2_0_1_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_2_0_1_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_2_0_1_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_2_0_1_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_2_0_1_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_2_0_1_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_2_0_1_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_2_0_1_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_2_0_1_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_2_0_1_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_2_0_1_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_2_0_1_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_0_2)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_2_0_2_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_2_0_2_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_2_0_2_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_2_0_2_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_2_0_2_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_2_0_2_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_2_0_2_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_2_0_2_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_2_0_2_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_2_0_2_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_2_0_2_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_2_0_2_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_2_0_2_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_2_0_2_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_2_0_2_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_2_0_2_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_2_0_2_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_2_0_2_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_2_0_2_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_2_0_2_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_2_0_2_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_2_0_2_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_2_0_2_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_2_0_2_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_2_0_2_string = "???????????";
    endcase
  end
  always @(*) begin
    case(LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size)
      MemAccessSize_B : LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size_string = "B";
      MemAccessSize_H : LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size_string = "H";
      MemAccessSize_W : LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size_string = "W";
      MemAccessSize_D : LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size_string = "D";
      default : LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_0_0)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_3_0_0_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_3_0_0_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_3_0_0_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_3_0_0_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_3_0_0_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_3_0_0_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_3_0_0_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_3_0_0_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_3_0_0_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_3_0_0_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_3_0_0_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_3_0_0_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_3_0_0_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_3_0_0_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_3_0_0_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_3_0_0_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_3_0_0_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_3_0_0_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_3_0_0_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_3_0_0_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_3_0_0_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_3_0_0_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_3_0_0_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_3_0_0_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_3_0_0_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_0_1)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_3_0_1_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_3_0_1_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_3_0_1_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_3_0_1_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_3_0_1_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_3_0_1_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_3_0_1_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_3_0_1_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_3_0_1_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_3_0_1_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_3_0_1_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_3_0_1_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_3_0_1_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_3_0_1_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_3_0_1_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_3_0_1_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_3_0_1_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_3_0_1_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_3_0_1_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_3_0_1_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_3_0_1_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_3_0_1_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_3_0_1_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_3_0_1_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_3_0_1_string = "???????????";
    endcase
  end
  always @(*) begin
    case(CommitPlugin_hw_robFlushPort_payload_reason)
      FlushReason_NONE : CommitPlugin_hw_robFlushPort_payload_reason_string = "NONE               ";
      FlushReason_FULL_FLUSH : CommitPlugin_hw_robFlushPort_payload_reason_string = "FULL_FLUSH         ";
      FlushReason_ROLLBACK_TO_ROB_IDX : CommitPlugin_hw_robFlushPort_payload_reason_string = "ROLLBACK_TO_ROB_IDX";
      default : CommitPlugin_hw_robFlushPort_payload_reason_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize)
      MemAccessSize_B : LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize_string = "B";
      MemAccessSize_H : LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize_string = "H";
      MemAccessSize_W : LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize_string = "W";
      MemAccessSize_D : LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize_string = "D";
      default : LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize)
      MemAccessSize_B : LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "B";
      MemAccessSize_H : LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "H";
      MemAccessSize_W : LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "W";
      MemAccessSize_D : LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "D";
      default : LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_hw_pushPortInst_payload_accessSize)
      MemAccessSize_B : StoreBufferPlugin_hw_pushPortInst_payload_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_hw_pushPortInst_payload_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_hw_pushPortInst_payload_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_hw_pushPortInst_payload_accessSize_string = "D";
      default : StoreBufferPlugin_hw_pushPortInst_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_hw_bypassQuerySizeIn)
      MemAccessSize_B : StoreBufferPlugin_hw_bypassQuerySizeIn_string = "B";
      MemAccessSize_H : StoreBufferPlugin_hw_bypassQuerySizeIn_string = "H";
      MemAccessSize_W : StoreBufferPlugin_hw_bypassQuerySizeIn_string = "W";
      MemAccessSize_D : StoreBufferPlugin_hw_bypassQuerySizeIn_string = "D";
      default : StoreBufferPlugin_hw_bypassQuerySizeIn_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size)
      MemAccessSize_B : StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size_string = "B";
      MemAccessSize_H : StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size_string = "H";
      MemAccessSize_W : StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size_string = "W";
      MemAccessSize_D : StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size_string = "D";
      default : StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size)
      MemAccessSize_B : LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size_string = "B";
      MemAccessSize_H : LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size_string = "H";
      MemAccessSize_W : LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size_string = "W";
      MemAccessSize_D : LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size_string = "D";
      default : LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size_string = "?";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_uopCode)
      BaseUopCode_NOP : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "MUL        ";
      BaseUopCode_DIV : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "IDLE       ";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit)
      ExeUnitType_NONE : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "FPU_DIV_SQRT       ";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_isa)
      IsaType_UNKNOWN : DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "UNKNOWN  ";
      IsaType_DEMO : DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "DEMO     ";
      IsaType_RISCV : DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "RISCV    ";
      IsaType_LOONGARCH : DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "LOONGARCH";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype)
      ArchRegType_GPR : DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "LA_CF";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype)
      ArchRegType_GPR : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "LA_CF";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype)
      ArchRegType_GPR : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "LA_CF";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_immUsage)
      ImmUsageType_NONE : DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "JUMP_OFFSET  ";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp)
      LogicOp_NONE : DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "XOR_1";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size)
      MemAccessSize_B : DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "B";
      MemAccessSize_H : DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "H";
      MemAccessSize_W : DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "W";
      MemAccessSize_D : DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "D";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition)
      BranchCondition_NUL : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LA_CF_FALSE";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "D";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "D";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest)
      MemAccessSize_B : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "D";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode)
      DecodeExCode_INVALID : DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "OK          ";
      default : DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode)
      BaseUopCode_NOP : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "MUL        ";
      BaseUopCode_DIV : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "IDLE       ";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit)
      ExeUnitType_NONE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "FPU_DIV_SQRT       ";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa)
      IsaType_UNKNOWN : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "UNKNOWN  ";
      IsaType_DEMO : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "DEMO     ";
      IsaType_RISCV : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "RISCV    ";
      IsaType_LOONGARCH : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "LOONGARCH";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype)
      ArchRegType_GPR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "LA_CF";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype)
      ArchRegType_GPR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "LA_CF";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype)
      ArchRegType_GPR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "LA_CF";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage)
      ImmUsageType_NONE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "JUMP_OFFSET  ";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp)
      LogicOp_NONE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "XOR_1";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size)
      MemAccessSize_B : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "B";
      MemAccessSize_H : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "H";
      MemAccessSize_W : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "W";
      MemAccessSize_D : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "D";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition)
      BranchCondition_NUL : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "LA_CF_FALSE";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "D";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "D";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest)
      MemAccessSize_B : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "D";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode)
      DecodeExCode_INVALID : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "OK          ";
      default : _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype)
      ArchRegType_GPR : DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype_string = "LA_CF";
      default : DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode)
      BaseUopCode_NOP : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "IDLE       ";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit)
      ExeUnitType_NONE : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_isa)
      IsaType_UNKNOWN : RobAllocPlugin_logic_allocatedUops_0_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : RobAllocPlugin_logic_allocatedUops_0_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : RobAllocPlugin_logic_allocatedUops_0_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : RobAllocPlugin_logic_allocatedUops_0_decoded_isa_string = "LOONGARCH";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype)
      ArchRegType_GPR : RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype_string = "LA_CF";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype)
      ArchRegType_GPR : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype_string = "LA_CF";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype)
      ArchRegType_GPR : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype_string = "LA_CF";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage)
      ImmUsageType_NONE : RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp)
      LogicOp_NONE : RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size)
      MemAccessSize_B : RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size_string = "D";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition)
      BranchCondition_NUL : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode_string = "OK          ";
      default : RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa)
      IsaType_UNKNOWN : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa_string = "LOONGARCH";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size_string = "D";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa)
      IsaType_UNKNOWN : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa_string = "LOONGARCH";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size_string = "D";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa)
      IsaType_UNKNOWN : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa_string = "LOONGARCH";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size_string = "D";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa)
      IsaType_UNKNOWN : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa_string = "LOONGARCH";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size_string = "D";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp)
      LogicOp_NONE : AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp_string = "XOR_1";
      default : AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage)
      ImmUsageType_NONE : AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string = "JUMP_OFFSET  ";
      default : AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa)
      IsaType_UNKNOWN : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa_string = "LOONGARCH";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size_string = "D";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition)
      BranchCondition_NUL : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "LA_CF_FALSE";
      default : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size)
      MemAccessSize_B : LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size_string = "B";
      MemAccessSize_H : LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size_string = "H";
      MemAccessSize_W : LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size_string = "W";
      MemAccessSize_D : LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size_string = "D";
      default : LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize)
      MemAccessSize_B : _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "B";
      MemAccessSize_H : _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "H";
      MemAccessSize_W : _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "W";
      MemAccessSize_D : _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "D";
      default : _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize)
      MemAccessSize_B : LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "B";
      MemAccessSize_H : LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "H";
      MemAccessSize_W : LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "W";
      MemAccessSize_D : LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "D";
      default : LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_combStage_payload_accessSize)
      MemAccessSize_B : io_outputs_0_combStage_payload_accessSize_string = "B";
      MemAccessSize_H : io_outputs_0_combStage_payload_accessSize_string = "H";
      MemAccessSize_W : io_outputs_0_combStage_payload_accessSize_string = "W";
      MemAccessSize_D : io_outputs_0_combStage_payload_accessSize_string = "D";
      default : io_outputs_0_combStage_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(io_outputs_1_combStage_payload_accessSize)
      MemAccessSize_B : io_outputs_1_combStage_payload_accessSize_string = "B";
      MemAccessSize_H : io_outputs_1_combStage_payload_accessSize_string = "H";
      MemAccessSize_W : io_outputs_1_combStage_payload_accessSize_string = "W";
      MemAccessSize_D : io_outputs_1_combStage_payload_accessSize_string = "D";
      default : io_outputs_1_combStage_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_outputs_0_combStage_translated_payload_size)
      MemAccessSize_B : _zz_io_outputs_0_combStage_translated_payload_size_string = "B";
      MemAccessSize_H : _zz_io_outputs_0_combStage_translated_payload_size_string = "H";
      MemAccessSize_W : _zz_io_outputs_0_combStage_translated_payload_size_string = "W";
      MemAccessSize_D : _zz_io_outputs_0_combStage_translated_payload_size_string = "D";
      default : _zz_io_outputs_0_combStage_translated_payload_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_combStage_translated_payload_size)
      MemAccessSize_B : io_outputs_0_combStage_translated_payload_size_string = "B";
      MemAccessSize_H : io_outputs_0_combStage_translated_payload_size_string = "H";
      MemAccessSize_W : io_outputs_0_combStage_translated_payload_size_string = "W";
      MemAccessSize_D : io_outputs_0_combStage_translated_payload_size_string = "D";
      default : io_outputs_0_combStage_translated_payload_size_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_outputs_1_combStage_translated_payload_accessSize)
      MemAccessSize_B : _zz_io_outputs_1_combStage_translated_payload_accessSize_string = "B";
      MemAccessSize_H : _zz_io_outputs_1_combStage_translated_payload_accessSize_string = "H";
      MemAccessSize_W : _zz_io_outputs_1_combStage_translated_payload_accessSize_string = "W";
      MemAccessSize_D : _zz_io_outputs_1_combStage_translated_payload_accessSize_string = "D";
      default : _zz_io_outputs_1_combStage_translated_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(io_outputs_1_combStage_translated_payload_accessSize)
      MemAccessSize_B : io_outputs_1_combStage_translated_payload_accessSize_string = "B";
      MemAccessSize_H : io_outputs_1_combStage_translated_payload_accessSize_string = "H";
      MemAccessSize_W : io_outputs_1_combStage_translated_payload_accessSize_string = "W";
      MemAccessSize_D : io_outputs_1_combStage_translated_payload_accessSize_string = "D";
      default : io_outputs_1_combStage_translated_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException)
      MemAccessSize_B : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_string = "B";
      MemAccessSize_H : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_string = "H";
      MemAccessSize_W : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_string = "W";
      MemAccessSize_D : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_string = "D";
      default : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize)
      MemAccessSize_B : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "B";
      MemAccessSize_H : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "H";
      MemAccessSize_W : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "W";
      MemAccessSize_D : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "D";
      default : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1)
      MemAccessSize_B : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1_string = "B";
      MemAccessSize_H : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1_string = "H";
      MemAccessSize_W : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1_string = "W";
      MemAccessSize_D : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1_string = "D";
      default : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2)
      MemAccessSize_B : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2_string = "B";
      MemAccessSize_H : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2_string = "H";
      MemAccessSize_W : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2_string = "W";
      MemAccessSize_D : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2_string = "D";
      default : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_pushCmd_payload_size)
      MemAccessSize_B : LoadQueuePlugin_logic_pushCmd_payload_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_pushCmd_payload_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_pushCmd_payload_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_pushCmd_payload_size_string = "D";
      default : LoadQueuePlugin_logic_pushCmd_payload_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slots_0_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slots_0_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slots_0_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slots_0_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slots_0_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slots_0_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slots_1_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slots_1_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slots_1_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slots_1_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slots_1_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slots_1_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slots_2_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slots_2_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slots_2_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slots_2_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slots_2_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slots_2_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slots_3_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slots_3_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slots_3_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slots_3_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slots_3_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slots_3_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slotsNext_0_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slotsNext_0_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slotsNext_0_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slotsNext_0_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slotsNext_0_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slotsNext_0_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slotsNext_1_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slotsNext_1_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slotsNext_1_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slotsNext_1_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slotsNext_1_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slotsNext_1_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slotsNext_2_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slotsNext_2_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slotsNext_2_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slotsNext_2_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slotsNext_2_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slotsNext_2_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_slotsNext_3_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_slotsNext_3_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_slotsNext_3_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_slotsNext_3_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_slotsNext_3_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_slotsNext_3_size_string = "?";
    endcase
  end
  always @(*) begin
    case(LoadQueuePlugin_logic_loadQueue_completingHead_size)
      MemAccessSize_B : LoadQueuePlugin_logic_loadQueue_completingHead_size_string = "B";
      MemAccessSize_H : LoadQueuePlugin_logic_loadQueue_completingHead_size_string = "H";
      MemAccessSize_W : LoadQueuePlugin_logic_loadQueue_completingHead_size_string = "W";
      MemAccessSize_D : LoadQueuePlugin_logic_loadQueue_completingHead_size_string = "D";
      default : LoadQueuePlugin_logic_loadQueue_completingHead_size_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slots_0_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slots_0_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slots_0_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slots_0_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slots_0_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slots_0_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slots_1_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slots_1_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slots_1_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slots_1_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slots_1_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slots_1_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slots_2_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slots_2_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slots_2_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slots_2_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slots_2_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slots_2_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slots_3_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slots_3_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slots_3_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slots_3_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slots_3_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slots_3_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slotsNext_0_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slotsNext_0_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slotsNext_0_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slotsNext_0_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slotsNext_0_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slotsNext_0_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slotsNext_1_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slotsNext_1_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slotsNext_1_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slotsNext_1_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slotsNext_1_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slotsNext_1_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slotsNext_2_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slotsNext_2_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slotsNext_2_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slotsNext_2_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slotsNext_2_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slotsNext_2_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(StoreBufferPlugin_logic_slotsNext_3_accessSize)
      MemAccessSize_B : StoreBufferPlugin_logic_slotsNext_3_accessSize_string = "B";
      MemAccessSize_H : StoreBufferPlugin_logic_slotsNext_3_accessSize_string = "H";
      MemAccessSize_W : StoreBufferPlugin_logic_slotsNext_3_accessSize_string = "W";
      MemAccessSize_D : StoreBufferPlugin_logic_slotsNext_3_accessSize_string = "D";
      default : StoreBufferPlugin_logic_slotsNext_3_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize)
      MemAccessSize_B : _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "B";
      MemAccessSize_H : _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "H";
      MemAccessSize_W : _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "W";
      MemAccessSize_D : _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "D";
      default : _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_ROBPlugin_aggregatedFlushSignal_payload_reason)
      FlushReason_NONE : _zz_ROBPlugin_aggregatedFlushSignal_payload_reason_string = "NONE               ";
      FlushReason_FULL_FLUSH : _zz_ROBPlugin_aggregatedFlushSignal_payload_reason_string = "FULL_FLUSH         ";
      FlushReason_ROLLBACK_TO_ROB_IDX : _zz_ROBPlugin_aggregatedFlushSignal_payload_reason_string = "ROLLBACK_TO_ROB_IDX";
      default : _zz_ROBPlugin_aggregatedFlushSignal_payload_reason_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(ICachePlugin_logic_refill_fsm_stateReg)
      ICachePlugin_logic_refill_fsm_BOOT : ICachePlugin_logic_refill_fsm_stateReg_string = "BOOT        ";
      ICachePlugin_logic_refill_fsm_IDLE : ICachePlugin_logic_refill_fsm_stateReg_string = "IDLE        ";
      ICachePlugin_logic_refill_fsm_SEND_REQ : ICachePlugin_logic_refill_fsm_stateReg_string = "SEND_REQ    ";
      ICachePlugin_logic_refill_fsm_RECEIVE_DATA : ICachePlugin_logic_refill_fsm_stateReg_string = "RECEIVE_DATA";
      ICachePlugin_logic_refill_fsm_COMMIT : ICachePlugin_logic_refill_fsm_stateReg_string = "COMMIT      ";
      default : ICachePlugin_logic_refill_fsm_stateReg_string = "????????????";
    endcase
  end
  always @(*) begin
    case(ICachePlugin_logic_refill_fsm_stateNext)
      ICachePlugin_logic_refill_fsm_BOOT : ICachePlugin_logic_refill_fsm_stateNext_string = "BOOT        ";
      ICachePlugin_logic_refill_fsm_IDLE : ICachePlugin_logic_refill_fsm_stateNext_string = "IDLE        ";
      ICachePlugin_logic_refill_fsm_SEND_REQ : ICachePlugin_logic_refill_fsm_stateNext_string = "SEND_REQ    ";
      ICachePlugin_logic_refill_fsm_RECEIVE_DATA : ICachePlugin_logic_refill_fsm_stateNext_string = "RECEIVE_DATA";
      ICachePlugin_logic_refill_fsm_COMMIT : ICachePlugin_logic_refill_fsm_stateNext_string = "COMMIT      ";
      default : ICachePlugin_logic_refill_fsm_stateNext_string = "????????????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    if(BpuPipelinePlugin_logic_u2_write_isFiring) begin
      if(BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken) begin
        _zz_1 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(BpuPipelinePlugin_logic_u2_write_isFiring) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
        if(when_ICachePlugin_l260_1) begin
          _zz_3 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_4 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
        if(when_ICachePlugin_l260) begin
          _zz_4 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_s1_PC_Gen_haltRequest_FetchPipelinePlugin2_l381 = 1'b0;
    if(when_FetchPipelinePlugin2_l380) begin
      _zz_s1_PC_Gen_haltRequest_FetchPipelinePlugin2_l381 = 1'b1;
    end
  end

  always @(*) begin
    when_Connection_l66 = 1'b0;
    if(FetchPipelinePlugin_doHardRedirect_listening) begin
      when_Connection_l66 = 1'b1;
    end
  end

  always @(*) begin
    _zz_s1_Rename_isFlushingRoot = 1'b0;
    if(FetchPipelinePlugin_doHardRedirect_listening) begin
      _zz_s1_Rename_isFlushingRoot = 1'b1;
    end
  end

  always @(*) begin
    _zz_s2_RobAlloc_haltRequest_RenamePlugin_l85 = 1'b0;
    if(when_RenamePlugin_l83) begin
      _zz_s2_RobAlloc_haltRequest_RenamePlugin_l85 = 1'b1;
    end
  end

  always @(*) begin
    _zz_s0_Decode_isFlushingRoot = 1'b0;
    if(FetchPipelinePlugin_doHardRedirect_listening) begin
      _zz_s0_Decode_isFlushingRoot = 1'b1;
    end
  end

  always @(*) begin
    CheckpointManagerPlugin_saveCheckpointTrigger = 1'b0;
    if(when_CommitPlugin_l216) begin
      CheckpointManagerPlugin_saveCheckpointTrigger = 1'b1;
    end
  end

  always @(*) begin
    CheckpointManagerPlugin_restoreCheckpointTrigger = 1'b0;
    if(when_CommitPlugin_l227) begin
      CheckpointManagerPlugin_restoreCheckpointTrigger = 1'b1;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_valid = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_valid = 1'b1;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_robPtr = 4'b0000;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_robPtr = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_robPtr;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx = 6'h0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_physDestIsFpr = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_physDestIsFpr = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_physDestIsFpr;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_writesToPhysReg = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_writesToPhysReg = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_writesToPhysReg;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_useSrc1 = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_useSrc1 = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_useSrc1;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_src1Data = 32'h0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_src1Data = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_src1Tag = 6'h0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_src1Tag = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Tag;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_src1Ready = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_src1Ready = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Ready;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_src1IsFpr = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_src1IsFpr = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1IsFpr;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_useSrc2 = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_useSrc2 = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_useSrc2;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_src2Data = 32'h0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_src2Data = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_src2Tag = 6'h0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_src2Tag = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Tag;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_src2Ready = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_src2Ready = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Ready;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_src2IsFpr = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_src2IsFpr = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2IsFpr;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_valid = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_valid = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_valid;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSub = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSub = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSub;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isAdd = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isAdd = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isAdd;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSigned = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSigned = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSigned;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp = LogicOp_NONE;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_valid = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_valid = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_valid;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRight = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRight = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRight;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isArithmetic = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isArithmetic = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isArithmetic;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRotate = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRotate = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRotate;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isDoubleWord = 1'b0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isDoubleWord = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isDoubleWord;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_imm = 32'h0;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_imm = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_imm;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_uop_immUsage = ImmUsageType_NONE;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_uop_immUsage = _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_data = _zz_AluIntEU_AluIntEuPlugin_euResult_data;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_writesToPreg = 1'bx;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_writesToPreg = _zz_AluIntEU_AluIntEuPlugin_euResult_writesToPreg;
    end
  end

  assign AluIntEU_AluIntEuPlugin_euResult_isMispredictedBranch = 1'bx;
  assign AluIntEU_AluIntEuPlugin_euResult_isTaken = 1'bx;
  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_hasException = 1'bx;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_hasException = _zz_AluIntEU_AluIntEuPlugin_euResult_hasException;
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_exceptionCode = 8'bxxxxxxxx;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_exceptionCode = {7'd0, _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_2};
    end
  end

  always @(*) begin
    AluIntEU_AluIntEuPlugin_euResult_destIsFpr = 1'bx;
    if(s3_Writeback_isFiring) begin
      AluIntEU_AluIntEuPlugin_euResult_destIsFpr = 1'b0;
    end
  end

  assign DispatchPlugin_logic_iqRegs_0_0_0 = BaseUopCode_ALU;
  assign DispatchPlugin_logic_iqRegs_0_0_1 = BaseUopCode_SHIFT;
  assign DispatchPlugin_logic_iqRegs_0_0_2 = BaseUopCode_NOP;
  assign DispatchPlugin_logic_iqRegs_0_0_3 = BaseUopCode_IDLE;
  always @(*) begin
    MulEU_MulEuPlugin_euResult_valid = 1'b0;
    if(mul_s7_Writeback_isFiring) begin
      MulEU_MulEuPlugin_euResult_valid = 1'b1;
    end
  end

  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_pc = 32'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_isValid = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_uopCode = BaseUopCode_NOP;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_exeUnit = ExeUnitType_NONE;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_isa = IsaType_UNKNOWN;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_idx = 5'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_archDest_rtype = ArchRegType_GPR;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_writeArchDestEn = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_idx = 5'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc1_rtype = ArchRegType_GPR;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_useArchSrc1 = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_idx = 5'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_archSrc2_rtype = ArchRegType_GPR;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_useArchSrc2 = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_usePcForAddr = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_imm = 32'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_immUsage = ImmUsageType_NONE;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_valid = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_isSub = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_isAdd = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_isSigned = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_aluCtrl_logicOp = LogicOp_NONE;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_valid = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_isRight = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_isArithmetic = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_isRotate = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_shiftCtrl_isDoubleWord = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_mulDivCtrl_valid = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_mulDivCtrl_isDiv = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_mulDivCtrl_isSigned = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_mulDivCtrl_isWordOp = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_size = MemAccessSize_W;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isSignedLoad = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isStore = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isLoadLinked = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isStoreCond = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_atomicOp = 5'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isFence = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_fenceMode = 8'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isCacheOp = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_cacheOpType = 5'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_memCtrl_isPrefetch = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_condition = BranchCondition_NUL;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_isJump = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_isLink = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_idx = 5'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_linkReg_rtype = ArchRegType_GPR;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_isIndirect = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchCtrl_laCfIdx = 3'b000;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_opType = 4'b0000;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc1 = MemAccessSize_W;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeSrc2 = MemAccessSize_W;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fpSizeDest = MemAccessSize_W;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_roundingMode = 3'b000;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_isIntegerDest = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_isSignedCvt = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fmaNegSrc1 = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_fpuCtrl_fcmpCond = 5'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_csrAddr = 14'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_isWrite = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_isRead = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_isExchange = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_csrCtrl_useUimmAsSrc = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_sysCtrl_sysCode = 20'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_sysCtrl_isExceptionReturn = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_sysCtrl_isTlbOp = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_sysCtrl_tlbOpType = 4'b0000;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_decodeExceptionCode = DecodeExCode_OK;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_hasDecodeException = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_isMicrocode = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_microcodeEntry = 8'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_isSerializing = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_isBranchOrJump = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchPrediction_isTaken = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchPrediction_target = 32'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_decoded_branchPrediction_wasPredicted = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_physSrc1_idx = 6'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_physSrc1IsFpr = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_physSrc2_idx = 6'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_physSrc2IsFpr = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_physDest_idx = 6'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_physDestIsFpr = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_oldPhysDest_idx = 6'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_oldPhysDestIsFpr = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_allocatesPhysDest = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_rename_writesToPhysReg = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_robPtr = 4'b0000;
  assign MulEU_MulEuPlugin_euResult_uop_uop_uniqueId = 16'h0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_dispatched = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_executed = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_hasException = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_uop_exceptionCode = 8'h0;
  always @(*) begin
    MulEU_MulEuPlugin_euResult_uop_robPtr = 4'b0000;
    if(mul_s7_Writeback_isFiring) begin
      MulEU_MulEuPlugin_euResult_uop_robPtr = _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_5;
    end
  end

  always @(*) begin
    MulEU_MulEuPlugin_euResult_uop_physDest_idx = 6'h0;
    if(mul_s7_Writeback_isFiring) begin
      MulEU_MulEuPlugin_euResult_uop_physDest_idx = _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_5;
    end
  end

  assign MulEU_MulEuPlugin_euResult_uop_physDestIsFpr = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_writesToPhysReg = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_useSrc1 = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_src1Data = 32'h0;
  assign MulEU_MulEuPlugin_euResult_uop_src1Tag = 6'h0;
  assign MulEU_MulEuPlugin_euResult_uop_src1Ready = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_src1IsFpr = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_useSrc2 = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_src2Data = 32'h0;
  assign MulEU_MulEuPlugin_euResult_uop_src2Tag = 6'h0;
  assign MulEU_MulEuPlugin_euResult_uop_src2Ready = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_src2IsFpr = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_mulDivCtrl_valid = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_mulDivCtrl_isDiv = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_mulDivCtrl_isSigned = 1'b0;
  assign MulEU_MulEuPlugin_euResult_uop_mulDivCtrl_isWordOp = 1'b0;
  always @(*) begin
    MulEU_MulEuPlugin_euResult_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(mul_s7_Writeback_isFiring) begin
      MulEU_MulEuPlugin_euResult_data = _zz_MulEU_MulEuPlugin_euResult_data_1[31:0];
    end
  end

  always @(*) begin
    MulEU_MulEuPlugin_euResult_writesToPreg = 1'bx;
    if(mul_s7_Writeback_isFiring) begin
      MulEU_MulEuPlugin_euResult_writesToPreg = _zz_MulEU_MulEuPlugin_euResult_writesToPreg_5;
    end
  end

  assign MulEU_MulEuPlugin_euResult_isMispredictedBranch = 1'bx;
  assign MulEU_MulEuPlugin_euResult_isTaken = 1'bx;
  always @(*) begin
    MulEU_MulEuPlugin_euResult_hasException = 1'bx;
    if(mul_s7_Writeback_isFiring) begin
      MulEU_MulEuPlugin_euResult_hasException = 1'b0;
    end
  end

  always @(*) begin
    MulEU_MulEuPlugin_euResult_exceptionCode = 8'bxxxxxxxx;
    if(mul_s7_Writeback_isFiring) begin
      MulEU_MulEuPlugin_euResult_exceptionCode = 8'h0;
    end
  end

  always @(*) begin
    MulEU_MulEuPlugin_euResult_destIsFpr = 1'bx;
    if(mul_s7_Writeback_isFiring) begin
      MulEU_MulEuPlugin_euResult_destIsFpr = 1'b0;
    end
  end

  assign DispatchPlugin_logic_iqRegs_1_0_0 = BaseUopCode_MUL;
  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_valid = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_valid = 1'b1;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_robPtr = 4'b0000;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_robPtr = _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_physDest_idx = 6'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_physDest_idx = _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr = _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg = _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_useSrc1 = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_useSrc1 = _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc1;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_src1Data = 32'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_src1Data = _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_src1Tag = 6'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_src1Tag = _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Tag;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_src1Ready = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_src1Ready = _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr = _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_useSrc2 = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_useSrc2 = _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc2;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_src2Data = 32'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_src2Data = _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_src2Tag = 6'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_src2Tag = _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Tag;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_src2Ready = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_src2Ready = _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr = _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition = BranchCondition_NUL;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx = 5'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype = ArchRegType_GPR;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx = 3'b000;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_imm = 32'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_imm = _zz_BranchEU_BranchEuPlugin_euResult_uop_imm;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_pc = 32'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_pc = _zz_BranchEU_BranchEuPlugin_euResult_uop_pc;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target = 32'h0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted = 1'b0;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted = _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_data = _zz_BranchEU_BranchEuPlugin_euResult_data;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_writesToPreg = 1'bx;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_writesToPreg = _zz_BranchEU_BranchEuPlugin_euResult_writesToPreg;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_isMispredictedBranch = 1'bx;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_isMispredictedBranch = _zz_BranchEU_BranchEuPlugin_euResult_isMispredictedBranch;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_isTaken = 1'bx;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_isTaken = _zz_BranchEU_BranchEuPlugin_euResult_isTaken;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_hasException = 1'bx;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_hasException = 1'b0;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_exceptionCode = 8'bxxxxxxxx;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_exceptionCode = 8'h0;
    end
  end

  always @(*) begin
    BranchEU_BranchEuPlugin_euResult_destIsFpr = 1'bx;
    if(s3_Result_isFiring) begin
      BranchEU_BranchEuPlugin_euResult_destIsFpr = 1'b0;
    end
  end

  assign DispatchPlugin_logic_iqRegs_2_0_0 = BaseUopCode_BRANCH;
  assign DispatchPlugin_logic_iqRegs_2_0_1 = BaseUopCode_JUMP_REG;
  assign DispatchPlugin_logic_iqRegs_2_0_2 = BaseUopCode_JUMP_IMM;
  always @(*) begin
    LsuEU_LsuEuPlugin_euResult_valid = 1'b0;
    if(when_LsuEuPlugin_l141) begin
      if(StoreBufferPlugin_hw_pushPortInst_fire) begin
        LsuEU_LsuEuPlugin_euResult_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    LsuEU_LsuEuPlugin_euResult_uop_robPtr = 4'b0000;
    if(when_LsuEuPlugin_l141) begin
      if(StoreBufferPlugin_hw_pushPortInst_fire) begin
        LsuEU_LsuEuPlugin_euResult_uop_robPtr = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr;
      end
    end
  end

  always @(*) begin
    LsuEU_LsuEuPlugin_euResult_uop_physDest_idx = 6'h0;
    if(when_LsuEuPlugin_l141) begin
      if(StoreBufferPlugin_hw_pushPortInst_fire) begin
        LsuEU_LsuEuPlugin_euResult_uop_physDest_idx = 6'h0;
      end
    end
  end

  assign LsuEU_LsuEuPlugin_euResult_uop_physDestIsFpr = 1'b0;
  always @(*) begin
    LsuEU_LsuEuPlugin_euResult_uop_writesToPhysReg = 1'b0;
    if(when_LsuEuPlugin_l141) begin
      if(StoreBufferPlugin_hw_pushPortInst_fire) begin
        LsuEU_LsuEuPlugin_euResult_uop_writesToPhysReg = 1'b0;
      end
    end
  end

  assign LsuEU_LsuEuPlugin_euResult_uop_useSrc1 = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_src1Data = 32'h0;
  assign LsuEU_LsuEuPlugin_euResult_uop_src1Tag = 6'h0;
  assign LsuEU_LsuEuPlugin_euResult_uop_src1Ready = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_src1IsFpr = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_useSrc2 = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_src2Data = 32'h0;
  assign LsuEU_LsuEuPlugin_euResult_uop_src2Tag = 6'h0;
  assign LsuEU_LsuEuPlugin_euResult_uop_src2Ready = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_src2IsFpr = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_size = MemAccessSize_W;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isSignedLoad = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isStore = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isLoadLinked = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isStoreCond = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_atomicOp = 5'h0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isFence = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_fenceMode = 8'h0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isCacheOp = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_cacheOpType = 5'h0;
  assign LsuEU_LsuEuPlugin_euResult_uop_memCtrl_isPrefetch = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_imm = 32'h0;
  assign LsuEU_LsuEuPlugin_euResult_uop_usePc = 1'b0;
  assign LsuEU_LsuEuPlugin_euResult_uop_pcData = 32'h0;
  assign LsuEU_LsuEuPlugin_euResult_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  always @(*) begin
    LsuEU_LsuEuPlugin_euResult_writesToPreg = 1'bx;
    if(when_LsuEuPlugin_l141) begin
      if(StoreBufferPlugin_hw_pushPortInst_fire) begin
        LsuEU_LsuEuPlugin_euResult_writesToPreg = 1'b0;
      end
    end
  end

  assign LsuEU_LsuEuPlugin_euResult_isMispredictedBranch = 1'bx;
  assign LsuEU_LsuEuPlugin_euResult_isTaken = 1'bx;
  always @(*) begin
    LsuEU_LsuEuPlugin_euResult_hasException = 1'bx;
    if(when_LsuEuPlugin_l141) begin
      if(StoreBufferPlugin_hw_pushPortInst_fire) begin
        LsuEU_LsuEuPlugin_euResult_hasException = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException;
      end
    end
  end

  always @(*) begin
    LsuEU_LsuEuPlugin_euResult_exceptionCode = 8'bxxxxxxxx;
    if(when_LsuEuPlugin_l141) begin
      if(StoreBufferPlugin_hw_pushPortInst_fire) begin
        LsuEU_LsuEuPlugin_euResult_exceptionCode = 8'h06;
      end
    end
  end

  always @(*) begin
    LsuEU_LsuEuPlugin_euResult_destIsFpr = 1'bx;
    if(when_LsuEuPlugin_l141) begin
      if(StoreBufferPlugin_hw_pushPortInst_fire) begin
        LsuEU_LsuEuPlugin_euResult_destIsFpr = 1'b0;
      end
    end
  end

  assign DispatchPlugin_logic_iqRegs_3_0_0 = BaseUopCode_LOAD;
  assign DispatchPlugin_logic_iqRegs_3_0_1 = BaseUopCode_STORE;
  assign DataCachePlugin_setup_writebackBusy = DataCachePlugin_setup_cache_io_writebackBusy;
  assign DataCachePlugin_setup_refillCompletions = DataCachePlugin_setup_cache_io_refillCompletions;
  always @(*) begin
    DataCachePlugin_setup_cache_io_mem_read_cmd_ready = io_mem_toAxi4_arCmdStaged_ready;
    if(when_Stream_l477) begin
      DataCachePlugin_setup_cache_io_mem_read_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! io_mem_toAxi4_arCmdStaged_valid);
  assign io_mem_toAxi4_arCmdStaged_valid = io_mem_read_cmd_rValid;
  assign io_mem_toAxi4_arCmdStaged_payload_id = io_mem_read_cmd_rData_id;
  assign io_mem_toAxi4_arCmdStaged_payload_address = io_mem_read_cmd_rData_address;
  assign DataCachePlugin_setup_dcacheMaster_ar_valid = io_mem_toAxi4_arCmdStaged_valid;
  assign DataCachePlugin_setup_dcacheMaster_ar_payload_addr = io_mem_toAxi4_arCmdStaged_payload_address;
  assign DataCachePlugin_setup_dcacheMaster_ar_payload_id = io_mem_toAxi4_arCmdStaged_payload_id;
  assign DataCachePlugin_setup_dcacheMaster_ar_payload_prot = 3'b010;
  assign DataCachePlugin_setup_dcacheMaster_ar_payload_len = 8'h07;
  assign DataCachePlugin_setup_dcacheMaster_ar_payload_size = 3'b010;
  assign DataCachePlugin_setup_dcacheMaster_ar_payload_burst = 2'b01;
  assign io_mem_toAxi4_arCmdStaged_ready = DataCachePlugin_setup_dcacheMaster_ar_ready;
  always @(*) begin
    DataCachePlugin_setup_dcacheMaster_r_ready = io_mem_toAxi4_rRspStaged_ready;
    if(when_Stream_l477_1) begin
      DataCachePlugin_setup_dcacheMaster_r_ready = 1'b1;
    end
  end

  assign when_Stream_l477_1 = (! io_mem_toAxi4_rRspStaged_valid);
  assign io_mem_toAxi4_rRspStaged_valid = DataCachePlugin_setup_dcacheMaster_r_rValid;
  assign io_mem_toAxi4_rRspStaged_payload_data = DataCachePlugin_setup_dcacheMaster_r_rData_data;
  assign io_mem_toAxi4_rRspStaged_payload_id = DataCachePlugin_setup_dcacheMaster_r_rData_id;
  assign io_mem_toAxi4_rRspStaged_payload_resp = DataCachePlugin_setup_dcacheMaster_r_rData_resp;
  assign io_mem_toAxi4_rRspStaged_payload_last = DataCachePlugin_setup_dcacheMaster_r_rData_last;
  assign DataCachePlugin_setup_cache_io_mem_read_rsp_payload_error = (! (io_mem_toAxi4_rRspStaged_payload_resp == 2'b00));
  assign io_mem_toAxi4_rRspStaged_ready = 1'b1;
  always @(*) begin
    DataCachePlugin_setup_cache_io_mem_write_cmd_ready = 1'b1;
    if(when_Stream_l1253) begin
      DataCachePlugin_setup_cache_io_mem_write_cmd_ready = 1'b0;
    end
    if(when_Stream_l1253_1) begin
      DataCachePlugin_setup_cache_io_mem_write_cmd_ready = 1'b0;
    end
  end

  assign when_Stream_l1253 = ((! io_mem_toAxi4_awRaw_ready) && io_mem_write_cmd_fork2_logic_linkEnable_0);
  assign when_Stream_l1253_1 = ((! io_mem_toAxi4_wRaw_ready) && io_mem_write_cmd_fork2_logic_linkEnable_1);
  assign io_mem_toAxi4_awRaw_valid = (DataCachePlugin_setup_cache_io_mem_write_cmd_valid && io_mem_write_cmd_fork2_logic_linkEnable_0);
  assign io_mem_toAxi4_awRaw_payload_last = DataCachePlugin_setup_cache_io_mem_write_cmd_payload_last;
  assign io_mem_toAxi4_awRaw_payload_fragment_address = DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_address;
  assign io_mem_toAxi4_awRaw_payload_fragment_data = DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_data;
  assign io_mem_toAxi4_awRaw_payload_fragment_id = DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_id;
  assign io_mem_toAxi4_awRaw_fire = (io_mem_toAxi4_awRaw_valid && io_mem_toAxi4_awRaw_ready);
  assign io_mem_toAxi4_wRaw_valid = (DataCachePlugin_setup_cache_io_mem_write_cmd_valid && io_mem_write_cmd_fork2_logic_linkEnable_1);
  assign io_mem_toAxi4_wRaw_payload_last = DataCachePlugin_setup_cache_io_mem_write_cmd_payload_last;
  assign io_mem_toAxi4_wRaw_payload_fragment_address = DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_address;
  assign io_mem_toAxi4_wRaw_payload_fragment_data = DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_data;
  assign io_mem_toAxi4_wRaw_payload_fragment_id = DataCachePlugin_setup_cache_io_mem_write_cmd_payload_fragment_id;
  assign io_mem_toAxi4_wRaw_fire = (io_mem_toAxi4_wRaw_valid && io_mem_toAxi4_wRaw_ready);
  assign when_Stream_l581 = (! io_mem_toAxi4_awRaw_payload_first);
  always @(*) begin
    io_mem_toAxi4_awFiltred_valid = io_mem_toAxi4_awRaw_valid;
    if(when_Stream_l581) begin
      io_mem_toAxi4_awFiltred_valid = 1'b0;
    end
  end

  always @(*) begin
    io_mem_toAxi4_awRaw_ready = io_mem_toAxi4_awFiltred_ready;
    if(when_Stream_l581) begin
      io_mem_toAxi4_awRaw_ready = 1'b1;
    end
  end

  assign io_mem_toAxi4_awFiltred_payload_last = io_mem_toAxi4_awRaw_payload_last;
  assign io_mem_toAxi4_awFiltred_payload_fragment_address = io_mem_toAxi4_awRaw_payload_fragment_address;
  assign io_mem_toAxi4_awFiltred_payload_fragment_data = io_mem_toAxi4_awRaw_payload_fragment_data;
  assign io_mem_toAxi4_awFiltred_payload_fragment_id = io_mem_toAxi4_awRaw_payload_fragment_id;
  always @(*) begin
    io_mem_toAxi4_awFiltred_ready = io_mem_toAxi4_aw_ready;
    if(when_Stream_l477_2) begin
      io_mem_toAxi4_awFiltred_ready = 1'b1;
    end
  end

  assign when_Stream_l477_2 = (! io_mem_toAxi4_aw_valid);
  assign io_mem_toAxi4_aw_valid = io_mem_toAxi4_awFiltred_rValid;
  assign io_mem_toAxi4_aw_payload_last = io_mem_toAxi4_awFiltred_rData_last;
  assign io_mem_toAxi4_aw_payload_fragment_address = io_mem_toAxi4_awFiltred_rData_fragment_address;
  assign io_mem_toAxi4_aw_payload_fragment_data = io_mem_toAxi4_awFiltred_rData_fragment_data;
  assign io_mem_toAxi4_aw_payload_fragment_id = io_mem_toAxi4_awFiltred_rData_fragment_id;
  assign DataCachePlugin_setup_dcacheMaster_aw_valid = io_mem_toAxi4_aw_valid;
  assign DataCachePlugin_setup_dcacheMaster_aw_payload_addr = io_mem_toAxi4_aw_payload_fragment_address;
  assign DataCachePlugin_setup_dcacheMaster_aw_payload_id = io_mem_toAxi4_aw_payload_fragment_id;
  assign DataCachePlugin_setup_dcacheMaster_aw_payload_prot = 3'b010;
  assign DataCachePlugin_setup_dcacheMaster_aw_payload_len = 8'h07;
  assign DataCachePlugin_setup_dcacheMaster_aw_payload_size = 3'b010;
  assign DataCachePlugin_setup_dcacheMaster_aw_payload_burst = 2'b01;
  assign io_mem_toAxi4_aw_ready = DataCachePlugin_setup_dcacheMaster_aw_ready;
  assign _zz_io_mem_toAxi4_wRaw_ready = (! io_mem_toAxi4_awFiltred_valid);
  assign io_mem_toAxi4_w_valid = (io_mem_toAxi4_wRaw_valid && _zz_io_mem_toAxi4_wRaw_ready);
  assign io_mem_toAxi4_wRaw_ready = (io_mem_toAxi4_w_ready && _zz_io_mem_toAxi4_wRaw_ready);
  assign io_mem_toAxi4_w_payload_last = io_mem_toAxi4_wRaw_payload_last;
  assign io_mem_toAxi4_w_payload_fragment_address = io_mem_toAxi4_wRaw_payload_fragment_address;
  assign io_mem_toAxi4_w_payload_fragment_data = io_mem_toAxi4_wRaw_payload_fragment_data;
  assign io_mem_toAxi4_w_payload_fragment_id = io_mem_toAxi4_wRaw_payload_fragment_id;
  always @(*) begin
    io_mem_toAxi4_w_ready = io_mem_toAxi4_wStaged_ready;
    if(when_Stream_l477_3) begin
      io_mem_toAxi4_w_ready = 1'b1;
    end
  end

  assign when_Stream_l477_3 = (! io_mem_toAxi4_wStaged_valid);
  assign io_mem_toAxi4_wStaged_valid = io_mem_toAxi4_w_rValid;
  assign io_mem_toAxi4_wStaged_payload_last = io_mem_toAxi4_w_rData_last;
  assign io_mem_toAxi4_wStaged_payload_fragment_address = io_mem_toAxi4_w_rData_fragment_address;
  assign io_mem_toAxi4_wStaged_payload_fragment_data = io_mem_toAxi4_w_rData_fragment_data;
  assign io_mem_toAxi4_wStaged_payload_fragment_id = io_mem_toAxi4_w_rData_fragment_id;
  assign DataCachePlugin_setup_dcacheMaster_w_valid = io_mem_toAxi4_wStaged_valid;
  assign DataCachePlugin_setup_dcacheMaster_w_payload_data = io_mem_toAxi4_wStaged_payload_fragment_data;
  assign DataCachePlugin_setup_dcacheMaster_w_payload_strb = 4'b1111;
  assign DataCachePlugin_setup_dcacheMaster_w_payload_last = io_mem_toAxi4_wStaged_payload_last;
  assign io_mem_toAxi4_wStaged_ready = DataCachePlugin_setup_dcacheMaster_w_ready;
  always @(*) begin
    DataCachePlugin_setup_dcacheMaster_b_ready = io_mem_toAxi4_bRspStaged_ready;
    if(when_Stream_l477_4) begin
      DataCachePlugin_setup_dcacheMaster_b_ready = 1'b1;
    end
  end

  assign when_Stream_l477_4 = (! io_mem_toAxi4_bRspStaged_valid);
  assign io_mem_toAxi4_bRspStaged_valid = DataCachePlugin_setup_dcacheMaster_b_rValid;
  assign io_mem_toAxi4_bRspStaged_payload_id = DataCachePlugin_setup_dcacheMaster_b_rData_id;
  assign io_mem_toAxi4_bRspStaged_payload_resp = DataCachePlugin_setup_dcacheMaster_b_rData_resp;
  assign DataCachePlugin_setup_cache_io_mem_write_rsp_payload_error = (! (io_mem_toAxi4_bRspStaged_payload_resp == 2'b00));
  assign io_mem_toAxi4_bRspStaged_ready = 1'b1;
  assign oneShot_13_io_triggerIn = (1'b1 && (_zz_when_Debug_l71 < _zz_io_triggerIn));
  assign _zz_when_Debug_l71_1 = 1'b1;
  assign when_Debug_l71 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_13);
  assign s0_Decode_isFiring = (s0_Decode_valid && s0_Decode_ready);
  assign oneShot_14_io_triggerIn = (s0_Decode_isFiring && (_zz_when_Debug_l71 < _zz_io_triggerIn_2));
  assign _zz_when_Debug_l71_2 = 5'h13;
  assign when_Debug_l71_1 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_1_1);
  assign s1_Rename_isFiring = (s1_Rename_valid && s1_Rename_ready);
  assign oneShot_15_io_triggerIn = (s1_Rename_isFiring && (_zz_when_Debug_l71 < _zz_io_triggerIn_4));
  assign _zz_when_Debug_l71_3 = 5'h15;
  assign when_Debug_l71_2 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_2_1);
  assign s2_RobAlloc_isFiring = (s2_RobAlloc_valid && s2_RobAlloc_ready);
  assign oneShot_16_io_triggerIn = (s2_RobAlloc_isFiring && (_zz_when_Debug_l71 < _zz_io_triggerIn_6));
  assign _zz_when_Debug_l71_4 = 5'h14;
  assign when_Debug_l71_3 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_3_1);
  assign s3_Dispatch_isFiring = (s3_Dispatch_valid && s3_Dispatch_ready);
  assign oneShot_17_io_triggerIn = (s3_Dispatch_isFiring && (_zz_when_Debug_l71 < _zz_io_triggerIn_8));
  assign _zz_when_Debug_l71_5 = 5'h16;
  assign when_Debug_l71_4 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_4_1);
  always @(*) begin
    CommitPlugin_hw_redirectPort_valid = 1'b0;
    if(when_CommitPlugin_l227) begin
      CommitPlugin_hw_redirectPort_valid = 1'b1;
    end
  end

  always @(*) begin
    CommitPlugin_hw_redirectPort_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_CommitPlugin_l227) begin
      CommitPlugin_hw_redirectPort_payload = ROBPlugin_robComponent_io_commit_0_entry_status_result;
    end
  end

  always @(*) begin
    BpuPipelinePlugin_updatePortIn_valid = 1'b0;
    if(when_CommitPlugin_l203) begin
      BpuPipelinePlugin_updatePortIn_valid = 1'b1;
    end
  end

  always @(*) begin
    BpuPipelinePlugin_updatePortIn_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_CommitPlugin_l203) begin
      BpuPipelinePlugin_updatePortIn_payload_pc = ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_pc;
    end
  end

  always @(*) begin
    BpuPipelinePlugin_updatePortIn_payload_isTaken = 1'bx;
    if(when_CommitPlugin_l203) begin
      BpuPipelinePlugin_updatePortIn_payload_isTaken = ROBPlugin_robComponent_io_commit_0_entry_status_isTaken;
    end
  end

  always @(*) begin
    BpuPipelinePlugin_updatePortIn_payload_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_CommitPlugin_l203) begin
      BpuPipelinePlugin_updatePortIn_payload_target = ROBPlugin_robComponent_io_commit_0_entry_status_result;
    end
  end

  assign CommitPlugin_maxCommitPcExt = 32'h80001000;
  assign CommitPlugin_maxCommitPcEnabledExt = 1'b1;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_valid = AluIntEU_AluIntEuPlugin_bypassOutputPort_valid;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_physRegIdx = AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_physRegIdx;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_physRegData = AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_physRegData;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_robPtr = AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_robPtr;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_isFPR = AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_isFPR;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_hasException = AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_hasException;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_payload_exceptionCode = AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_exceptionCode;
  assign MulEU_MulEuPlugin_bypassOutputPort_toStream_valid = MulEU_MulEuPlugin_bypassOutputPort_valid;
  assign MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_physRegIdx = MulEU_MulEuPlugin_bypassOutputPort_payload_physRegIdx;
  assign MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_physRegData = MulEU_MulEuPlugin_bypassOutputPort_payload_physRegData;
  assign MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_robPtr = MulEU_MulEuPlugin_bypassOutputPort_payload_robPtr;
  assign MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_isFPR = MulEU_MulEuPlugin_bypassOutputPort_payload_isFPR;
  assign MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_hasException = MulEU_MulEuPlugin_bypassOutputPort_payload_hasException;
  assign MulEU_MulEuPlugin_bypassOutputPort_toStream_payload_exceptionCode = MulEU_MulEuPlugin_bypassOutputPort_payload_exceptionCode;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_toStream_valid = BranchEU_BranchEuPlugin_bypassOutputPort_valid;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_physRegIdx = BranchEU_BranchEuPlugin_bypassOutputPort_payload_physRegIdx;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_physRegData = BranchEU_BranchEuPlugin_bypassOutputPort_payload_physRegData;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_robPtr = BranchEU_BranchEuPlugin_bypassOutputPort_payload_robPtr;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_isFPR = BranchEU_BranchEuPlugin_bypassOutputPort_payload_isFPR;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_hasException = BranchEU_BranchEuPlugin_bypassOutputPort_payload_hasException;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_toStream_payload_exceptionCode = BranchEU_BranchEuPlugin_bypassOutputPort_payload_exceptionCode;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_toStream_ready = streamArbiter_8_io_inputs_0_ready;
  assign MulEU_MulEuPlugin_bypassOutputPort_toStream_ready = streamArbiter_8_io_inputs_1_ready;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_toStream_ready = streamArbiter_8_io_inputs_2_ready;
  assign io_output_combStage_valid = streamArbiter_8_io_output_valid;
  assign io_output_combStage_payload_physRegIdx = streamArbiter_8_io_output_payload_physRegIdx;
  assign io_output_combStage_payload_physRegData = streamArbiter_8_io_output_payload_physRegData;
  assign io_output_combStage_payload_robPtr = streamArbiter_8_io_output_payload_robPtr;
  assign io_output_combStage_payload_isFPR = streamArbiter_8_io_output_payload_isFPR;
  assign io_output_combStage_payload_hasException = streamArbiter_8_io_output_payload_hasException;
  assign io_output_combStage_payload_exceptionCode = streamArbiter_8_io_output_payload_exceptionCode;
  assign io_output_combStage_ready = 1'b1;
  assign AguPlugin_logic_bypassFlow_valid = io_output_combStage_valid;
  assign AguPlugin_logic_bypassFlow_payload_physRegIdx = io_output_combStage_payload_physRegIdx;
  assign AguPlugin_logic_bypassFlow_payload_physRegData = io_output_combStage_payload_physRegData;
  assign AguPlugin_logic_bypassFlow_payload_robPtr = io_output_combStage_payload_robPtr;
  assign AguPlugin_logic_bypassFlow_payload_isFPR = io_output_combStage_payload_isFPR;
  assign AguPlugin_logic_bypassFlow_payload_hasException = io_output_combStage_payload_hasException;
  assign AguPlugin_logic_bypassFlow_payload_exceptionCode = io_output_combStage_payload_exceptionCode;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_0 = 6'h0;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_1 = 6'h01;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_2 = 6'h02;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_3 = 6'h03;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_4 = 6'h04;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_5 = 6'h05;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_6 = 6'h06;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_7 = 6'h07;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_8 = 6'h08;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_9 = 6'h09;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_10 = 6'h0a;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_11 = 6'h0b;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_12 = 6'h0c;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_13 = 6'h0d;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_14 = 6'h0e;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_15 = 6'h0f;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_16 = 6'h10;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_17 = 6'h11;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_18 = 6'h12;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_19 = 6'h13;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_20 = 6'h14;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_21 = 6'h15;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_22 = 6'h16;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_23 = 6'h17;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_24 = 6'h18;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_25 = 6'h19;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_26 = 6'h1a;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_27 = 6'h1b;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_28 = 6'h1c;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_29 = 6'h1d;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_30 = 6'h1e;
  assign CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_31 = 6'h1f;
  assign _zz_220 = zz_CheckpointManagerPlugin_logic_initialFreeMask(1'b0);
  always @(*) CheckpointManagerPlugin_logic_initialFreeMask = _zz_220;
  assign CheckpointManagerPlugin_logic_initialBtCheckpoint_busyBits = 64'h0;
  always @(*) begin
    CommitPlugin_hw_robFlushPort_valid = 1'b0;
    if(when_CommitPlugin_l227) begin
      CommitPlugin_hw_robFlushPort_valid = 1'b1;
    end
  end

  always @(*) begin
    CommitPlugin_hw_robFlushPort_payload_reason = (2'bxx);
    if(when_CommitPlugin_l227) begin
      CommitPlugin_hw_robFlushPort_payload_reason = FlushReason_FULL_FLUSH;
    end
  end

  always @(*) begin
    CommitPlugin_hw_robFlushPort_payload_targetRobPtr = 4'bxxxx;
    if(when_CommitPlugin_l227) begin
      CommitPlugin_hw_robFlushPort_payload_targetRobPtr = 4'bxxxx;
    end
  end

  always @(*) begin
    CommitPlugin_hw_busyTableClearPort_valid = 1'b0;
    if(when_CommitPlugin_l265) begin
      CommitPlugin_hw_busyTableClearPort_valid = 1'b1;
    end
  end

  always @(*) begin
    CommitPlugin_hw_busyTableClearPort_payload = 6'bxxxxxx;
    if(when_CommitPlugin_l265) begin
      CommitPlugin_hw_busyTableClearPort_payload = ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_oldPhysDest_idx;
    end
  end

  assign CommitPlugin_logic_s0_isMispredictedBranch = ((((CommitPlugin_commitEnableExt && ROBPlugin_robComponent_io_commit_0_valid) && ROBPlugin_robComponent_io_commit_0_entry_status_done) && ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isBranchOrJump) && ROBPlugin_robComponent_io_commit_0_entry_status_isMispredictedBranch);
  always @(*) begin
    CommitPlugin_logic_s0_commitAckMasks_0 = 1'b0;
    if(when_CommitPlugin_l216) begin
      CommitPlugin_logic_s0_commitAckMasks_0 = 1'b1;
    end
    if(when_CommitPlugin_l227) begin
      CommitPlugin_logic_s0_commitAckMasks_0 = 1'b0;
    end
  end

  assign when_CommitPlugin_l203 = (((CommitPlugin_commitEnableExt && ROBPlugin_robComponent_io_commit_0_valid) && ROBPlugin_robComponent_io_commit_0_entry_status_done) && ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isBranchOrJump);
  assign when_CommitPlugin_l216 = (((CommitPlugin_commitEnableExt && ROBPlugin_robComponent_io_commit_0_valid) && ROBPlugin_robComponent_io_commit_0_entry_status_done) && (! CommitPlugin_logic_s0_isMispredictedBranch));
  assign when_CommitPlugin_l227 = (((CommitPlugin_commitEnableExt && ROBPlugin_robComponent_io_commit_0_valid) && ROBPlugin_robComponent_io_commit_0_entry_status_done) && CommitPlugin_logic_s0_isMispredictedBranch);
  assign when_CommitPlugin_l265 = (CommitPlugin_logic_s0_commitAckMasks_0 && ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_allocatesPhysDest);
  assign CommitPlugin_logic_s0_committedThisCycle_comb = _zz_CommitPlugin_logic_s0_committedThisCycle_comb;
  assign CommitPlugin_logic_s0_recycledThisCycle_comb = _zz_CommitPlugin_logic_s0_recycledThisCycle_comb;
  assign CommitPlugin_logic_s0_flushedThisCycle_comb = CommitPlugin_hw_robFlushPort_valid;
  assign CommitPlugin_logic_s0_commitPcs_0 = ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_pc;
  assign CommitPlugin_logic_s0_maxCommitPcThisCycle = (CommitPlugin_logic_s0_commitAckMasks_0 ? CommitPlugin_logic_s0_commitPcs_0 : 32'h0);
  assign CommitPlugin_logic_s0_anyCommitOOB = (CommitPlugin_maxCommitPcEnabledExt && (CommitPlugin_logic_s0_commitAckMasks_0 && (CommitPlugin_maxCommitPcExt < CommitPlugin_logic_s0_commitPcs_0)));
  assign CommitPlugin_logic_s0_commitSlotLogs_0_valid = ROBPlugin_robComponent_io_commit_0_valid;
  assign CommitPlugin_logic_s0_commitSlotLogs_0_canCommit = (ROBPlugin_robComponent_io_commit_0_canCommit && CommitPlugin_commitEnableExt);
  assign CommitPlugin_logic_s0_commitSlotLogs_0_doCommit = CommitPlugin_logic_s0_commitAckMasks_0;
  assign CommitPlugin_logic_s0_commitSlotLogs_0_robPtr = ROBPlugin_robComponent_io_commit_0_entry_payload_uop_robPtr;
  assign CommitPlugin_logic_s0_commitSlotLogs_0_oldPhysDest = ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_oldPhysDest_idx;
  assign CommitPlugin_logic_s0_commitSlotLogs_0_allocatesPhysDest = ROBPlugin_robComponent_io_commit_0_entry_payload_uop_rename_allocatesPhysDest;
  assign CommitPlugin_logic_s1_s1_hasCommitsThisCycle = (1'b0 < CommitPlugin_logic_s1_s1_committedThisCycle);
  assign when_CommitPlugin_l317 = (CommitPlugin_logic_s1_s1_hasCommitsThisCycle && (CommitPlugin_maxCommitPcReg < CommitPlugin_logic_s1_s1_maxCommitPcThisCycle));
  assign oneShot_18_io_triggerIn = (CommitPlugin_logic_s0_committedThisCycle_comb[0] && (_zz_when_Debug_l71 < _zz_io_triggerIn_10));
  assign _zz_when_Debug_l71_6 = 5'h19;
  assign when_Debug_l71_5 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_5_1);
  assign _zz_26 = 8'he3;
  assign lA32RSimpleDecoder_1_io_pcIn = (s0_Decode_IssuePipelineSignals_GROUP_PC_IN + 32'h0);
  always @(*) begin
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isValid = lA32RSimpleDecoder_1_io_decodedUop_isValid;
    if(when_DecodePlugin_l66) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isValid = 1'b0;
    end
    if(s0_Decode_IssuePipelineSignals_IS_FAULT_IN) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isValid = 1'b0;
    end
    if(when_DecodePlugin_l79) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isValid = 1'b0;
    end
  end

  always @(*) begin
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode = lA32RSimpleDecoder_1_io_decodedUop_uopCode;
    if(s0_Decode_IssuePipelineSignals_IS_FAULT_IN) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode = BaseUopCode_ILLEGAL;
    end
  end

  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit = lA32RSimpleDecoder_1_io_decodedUop_exeUnit;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa = lA32RSimpleDecoder_1_io_decodedUop_isa;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype = lA32RSimpleDecoder_1_io_decodedUop_archDest_rtype;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_writeArchDestEn = lA32RSimpleDecoder_1_io_decodedUop_writeArchDestEn;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype = lA32RSimpleDecoder_1_io_decodedUop_archSrc1_rtype;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_idx = lA32RSimpleDecoder_1_io_decodedUop_archSrc2_idx;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype = lA32RSimpleDecoder_1_io_decodedUop_archSrc2_rtype;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage = lA32RSimpleDecoder_1_io_decodedUop_immUsage;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp = lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_logicOp;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_size;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition = lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_condition;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype = lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_linkReg_rtype;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1 = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeSrc1;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2 = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeSrc2;
  assign _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fpSizeDest;
  always @(*) begin
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode = lA32RSimpleDecoder_1_io_decodedUop_decodeExceptionCode;
    if(s0_Decode_IssuePipelineSignals_IS_FAULT_IN) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode = DecodeExCode_FETCH_ERROR;
    end
  end

  always @(*) begin
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_hasDecodeException = lA32RSimpleDecoder_1_io_decodedUop_hasDecodeException;
    if(s0_Decode_IssuePipelineSignals_IS_FAULT_IN) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_hasDecodeException = 1'b1;
    end
  end

  always @(*) begin
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken = lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_isTaken;
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken = 1'bx;
    if(when_DecodePlugin_l85) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken = s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_isTaken;
    end
  end

  always @(*) begin
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target = lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_target;
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_DecodePlugin_l85) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target = s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_target;
    end
  end

  always @(*) begin
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted = lA32RSimpleDecoder_1_io_decodedUop_branchPrediction_wasPredicted;
    _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted = 1'bx;
    if(when_DecodePlugin_l85) begin
      _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted = s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_wasPredicted;
    end
  end

  assign when_DecodePlugin_l66 = ((((_zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode == BaseUopCode_ALU) || (_zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode == BaseUopCode_SHIFT)) && (! _zz_DecodePlugin_logic_decodedUopsOutputVec_0_writeArchDestEn)) || (_zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode == BaseUopCode_NOP));
  assign when_DecodePlugin_l79 = (! s0_Decode_IssuePipelineSignals_VALID_MASK[0]);
  assign when_DecodePlugin_l85 = (! when_DecodePlugin_l66);
  assign DecodePlugin_logic_decodedUopsOutputVec_0_pc = lA32RSimpleDecoder_1_io_decodedUop_pc;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_isValid = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isValid;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_uopCode = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_uopCode;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_isa = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_isa;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_archDest_idx = lA32RSimpleDecoder_1_io_decodedUop_archDest_idx;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_writeArchDestEn = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_writeArchDestEn;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_idx = lA32RSimpleDecoder_1_io_decodedUop_archSrc1_idx;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_useArchSrc1 = lA32RSimpleDecoder_1_io_decodedUop_useArchSrc1;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_idx = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_idx;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_useArchSrc2 = lA32RSimpleDecoder_1_io_decodedUop_useArchSrc2;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_usePcForAddr = lA32RSimpleDecoder_1_io_decodedUop_usePcForAddr;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_imm = lA32RSimpleDecoder_1_io_decodedUop_imm;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_immUsage = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_immUsage;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_valid = lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_valid;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isSub = lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isSub;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isAdd = lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isAdd;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isSigned = lA32RSimpleDecoder_1_io_decodedUop_aluCtrl_isSigned;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_valid = lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_valid;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isRight = lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isRight;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isArithmetic = lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isArithmetic;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isRotate = lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isRotate;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isDoubleWord = lA32RSimpleDecoder_1_io_decodedUop_shiftCtrl_isDoubleWord;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_valid = lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_valid;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isDiv = lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isDiv;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isSigned = lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isSigned;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isWordOp = lA32RSimpleDecoder_1_io_decodedUop_mulDivCtrl_isWordOp;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isSignedLoad = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isSignedLoad;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isStore = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isStore;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isLoadLinked = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isLoadLinked;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isStoreCond = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isStoreCond;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_atomicOp = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_atomicOp;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isFence = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isFence;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_fenceMode = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_fenceMode;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isCacheOp = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isCacheOp;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_cacheOpType = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_cacheOpType;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isPrefetch = lA32RSimpleDecoder_1_io_decodedUop_memCtrl_isPrefetch;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isJump = lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isJump;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isLink = lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isLink;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_idx = lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_linkReg_idx;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isIndirect = lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_isIndirect;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_laCfIdx = lA32RSimpleDecoder_1_io_decodedUop_branchCtrl_laCfIdx;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_opType = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_opType;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1 = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2 = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_roundingMode = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_roundingMode;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_isIntegerDest = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_isIntegerDest;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_isSignedCvt = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_isSignedCvt;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fmaNegSrc1 = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fmaNegSrc1;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fcmpCond = lA32RSimpleDecoder_1_io_decodedUop_fpuCtrl_fcmpCond;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_csrAddr = lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_csrAddr;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isWrite = lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isWrite;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isRead = lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isRead;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isExchange = lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_isExchange;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_useUimmAsSrc = lA32RSimpleDecoder_1_io_decodedUop_csrCtrl_useUimmAsSrc;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_sysCode = lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_sysCode;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_isExceptionReturn = lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_isExceptionReturn;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_isTlbOp = lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_isTlbOp;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_tlbOpType = lA32RSimpleDecoder_1_io_decodedUop_sysCtrl_tlbOpType;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_hasDecodeException = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_hasDecodeException;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_isMicrocode = lA32RSimpleDecoder_1_io_decodedUop_isMicrocode;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_microcodeEntry = lA32RSimpleDecoder_1_io_decodedUop_microcodeEntry;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_isSerializing = lA32RSimpleDecoder_1_io_decodedUop_isSerializing;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_isBranchOrJump = lA32RSimpleDecoder_1_io_decodedUop_isBranchOrJump;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target;
  assign DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted = _zz_DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_pc = DecodePlugin_logic_decodedUopsOutputVec_0_pc;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isValid = DecodePlugin_logic_decodedUopsOutputVec_0_isValid;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode = DecodePlugin_logic_decodedUopsOutputVec_0_uopCode;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit = DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa = DecodePlugin_logic_decodedUopsOutputVec_0_isa;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx = DecodePlugin_logic_decodedUopsOutputVec_0_archDest_idx;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype = DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn = DecodePlugin_logic_decodedUopsOutputVec_0_writeArchDestEn;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx = DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_idx;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype = DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1 = DecodePlugin_logic_decodedUopsOutputVec_0_useArchSrc1;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx = DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_idx;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype = DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2 = DecodePlugin_logic_decodedUopsOutputVec_0_useArchSrc2;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr = DecodePlugin_logic_decodedUopsOutputVec_0_usePcForAddr;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_imm = DecodePlugin_logic_decodedUopsOutputVec_0_imm;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage = DecodePlugin_logic_decodedUopsOutputVec_0_immUsage;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid = DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_valid;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub = DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isSub;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd = DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isAdd;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned = DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isSigned;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp = DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid = DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_valid;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight = DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isRight;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic = DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isArithmetic;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate = DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isRotate;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord = DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isDoubleWord;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid = DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_valid;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv = DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isDiv;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned = DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isSigned;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp = DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isWordOp;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isSignedLoad;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isStore;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isLoadLinked;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isStoreCond;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_atomicOp;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isFence;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_fenceMode;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isCacheOp;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_cacheOpType;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch = DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isPrefetch;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition = DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump = DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isJump;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink = DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isLink;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx = DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_idx;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype = DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect = DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isIndirect;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx = DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_laCfIdx;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_opType;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1 = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2 = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_roundingMode;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_isIntegerDest;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_isSignedCvt;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1 = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fmaNegSrc1;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond = DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fcmpCond;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr = DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_csrAddr;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite = DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isWrite;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead = DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isRead;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange = DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isExchange;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc = DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_useUimmAsSrc;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode = DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_sysCode;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn = DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_isExceptionReturn;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp = DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_isTlbOp;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType = DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_tlbOpType;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode = DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException = DecodePlugin_logic_decodedUopsOutputVec_0_hasDecodeException;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode = DecodePlugin_logic_decodedUopsOutputVec_0_isMicrocode;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry = DecodePlugin_logic_decodedUopsOutputVec_0_microcodeEntry;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isSerializing = DecodePlugin_logic_decodedUopsOutputVec_0_isSerializing;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump = DecodePlugin_logic_decodedUopsOutputVec_0_isBranchOrJump;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken = DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target = DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target;
  assign s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted = DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted;
  assign when_DecodePlugin_l117 = (s0_Decode_isFiring && DecodePlugin_logic_decodedUopsOutputVec_0_isValid);
  assign _zz_27 = (DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype == ArchRegType_GPR);
  assign _zz_28 = (DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype == ArchRegType_FPR);
  assign _zz_29 = (DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype == ArchRegType_CSR);
  assign _zz_30 = (DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype == ArchRegType_GPR);
  assign _zz_31 = (DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype == ArchRegType_FPR);
  assign _zz_32 = (DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype == ArchRegType_CSR);
  assign _zz_33 = (DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype == ArchRegType_GPR);
  assign _zz_34 = (DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype == ArchRegType_FPR);
  assign _zz_35 = (DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype == ArchRegType_CSR);
  assign _zz_36 = (DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype == ArchRegType_GPR);
  assign _zz_37 = (DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype == ArchRegType_FPR);
  assign _zz_38 = (DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype == ArchRegType_CSR);
  assign SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_enable = (s1_Rename_valid && s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn);
  assign s1_Rename_IssuePipelineSignals_NEEDS_PHYS_REG_0 = s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn;
  assign RenamePlugin_logic_s2_logic_allocationOk = (&((! s2_RobAlloc_IssuePipelineSignals_NEEDS_PHYS_REG_0) || SimpleFreeListPlugin_early_setup_freeList_io_allocate_0_success));
  assign when_RenamePlugin_l83 = (s2_RobAlloc_valid && (! RenamePlugin_logic_s2_logic_allocationOk));
  assign _zz_39 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype == ArchRegType_GPR);
  assign _zz_40 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype == ArchRegType_FPR);
  assign _zz_41 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype == ArchRegType_CSR);
  assign _zz_42 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype == ArchRegType_GPR);
  assign _zz_43 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype == ArchRegType_FPR);
  assign _zz_44 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype == ArchRegType_CSR);
  assign _zz_45 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype == ArchRegType_GPR);
  assign _zz_46 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype == ArchRegType_FPR);
  assign _zz_47 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype == ArchRegType_CSR);
  assign _zz_48 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype == ArchRegType_GPR);
  assign _zz_49 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype == ArchRegType_FPR);
  assign _zz_50 = (s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype == ArchRegType_CSR);
  assign s2_RobAlloc_haltRequest_RenamePlugin_l85 = _zz_s2_RobAlloc_haltRequest_RenamePlugin_l85;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_pc = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_pc;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isValid = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isValid;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_uopCode;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_exeUnit;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isa;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_idx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archDest_idx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archDest_rtype;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_writeArchDestEn = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_writeArchDestEn;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_idx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc1_idx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc1_rtype;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_useArchSrc1 = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_useArchSrc1;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_idx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc2_idx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_archSrc2_rtype;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_useArchSrc2 = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_useArchSrc2;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_usePcForAddr = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_usePcForAddr;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_imm = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_imm;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_immUsage;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_valid = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_valid;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isSub = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isSub;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isAdd = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isAdd;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isSigned = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_isSigned;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_aluCtrl_logicOp;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_valid = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_valid;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isRight = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isRight;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isArithmetic = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isArithmetic;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isRotate = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isRotate;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isDoubleWord = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_shiftCtrl_isDoubleWord;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_valid = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_valid;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isDiv = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isDiv;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isSigned = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isSigned;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isWordOp = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_mulDivCtrl_isWordOp;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_size;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isSignedLoad = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isSignedLoad;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isStore = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isStore;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isLoadLinked = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isLoadLinked;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isStoreCond = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isStoreCond;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_atomicOp = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_atomicOp;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isFence = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isFence;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_fenceMode = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_fenceMode;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isCacheOp = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isCacheOp;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_cacheOpType = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_cacheOpType;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isPrefetch = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_memCtrl_isPrefetch;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_condition;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isJump = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isJump;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isLink = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isLink;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_idx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_linkReg_idx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isIndirect = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_isIndirect;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_laCfIdx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchCtrl_laCfIdx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_opType = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_opType;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1 = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2 = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_roundingMode = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_roundingMode;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_isIntegerDest = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_isIntegerDest;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_isSignedCvt = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_isSignedCvt;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1 = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fmaNegSrc1;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fcmpCond = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_fpuCtrl_fcmpCond;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_csrAddr = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_csrAddr;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isWrite = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isWrite;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isRead = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isRead;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isExchange = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_isExchange;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_useUimmAsSrc = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_csrCtrl_useUimmAsSrc;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_sysCode = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_sysCode;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_isExceptionReturn = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_isExceptionReturn;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_isTlbOp = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_isTlbOp;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_tlbOpType = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_sysCtrl_tlbOpType;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_decodeExceptionCode;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_hasDecodeException = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_hasDecodeException;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isMicrocode = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isMicrocode;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_microcodeEntry = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_microcodeEntry;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isSerializing = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isSerializing;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isBranchOrJump = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_isBranchOrJump;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_isTaken = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_isTaken;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_target = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_target;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_wasPredicted = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_decoded_branchPrediction_wasPredicted;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc1_idx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc1_idx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc1IsFpr = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc1IsFpr;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc2_idx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc2_idx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc2IsFpr = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physSrc2IsFpr;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physDest_idx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physDest_idx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physDestIsFpr = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physDestIsFpr;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_oldPhysDest_idx = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_oldPhysDest_idx;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_oldPhysDestIsFpr = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_oldPhysDestIsFpr;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_allocatesPhysDest = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_allocatesPhysDest;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_writesToPhysReg = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_writesToPhysReg;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_robPtr = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_robPtr;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_uniqueId = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_uniqueId;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_dispatched = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_dispatched;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_executed = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_executed;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_hasException = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_hasException;
  assign s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_exceptionCode = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_exceptionCode;
  assign RenameMapTablePlugin_early_setup_rat_io_writePorts_0_wen = (s2_RobAlloc_isFiring && RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_allocatesPhysDest);
  assign RenamePlugin_setup_btSetBusyPorts_0_valid = (s2_RobAlloc_isFiring && RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_allocatesPhysDest);
  assign RenamePlugin_setup_btSetBusyPorts_0_payload = RenamePlugin_setup_renameUnit_io_renamedUopsOut_0_rename_physDest_idx;
  assign s2_RobAlloc_haltRequest_RobAllocPlugin_l30 = (! ROBPlugin_robComponent_io_allocate_0_ready);
  assign ROBPlugin_robComponent_io_allocate_0_valid = (s2_RobAlloc_isFiring && s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isValid);
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_pc = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_pc;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_isValid = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isValid;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_uopCode;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_exeUnit;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_isa = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isa;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_idx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_idx;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archDest_rtype;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_writeArchDestEn = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_writeArchDestEn;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_idx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_idx;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc1_rtype;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_useArchSrc1 = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_useArchSrc1;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_idx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_idx;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_archSrc2_rtype;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_useArchSrc2 = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_useArchSrc2;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_usePcForAddr = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_usePcForAddr;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_imm = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_imm;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_immUsage;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_valid = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_valid;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isSub = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isSub;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isAdd = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isAdd;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isSigned = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_isSigned;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_aluCtrl_logicOp;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_valid = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_valid;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isRight = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isRight;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isArithmetic = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isArithmetic;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isRotate = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isRotate;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isDoubleWord = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_valid = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_valid;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isDiv = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isDiv;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isSigned = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isSigned;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isWordOp = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_mulDivCtrl_isWordOp;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_size;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isSignedLoad = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isSignedLoad;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isStore = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isStore;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isLoadLinked = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isLoadLinked;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isStoreCond = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isStoreCond;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_atomicOp = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_atomicOp;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isFence = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isFence;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_fenceMode = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_fenceMode;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isCacheOp = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isCacheOp;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_cacheOpType = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_cacheOpType;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isPrefetch = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_memCtrl_isPrefetch;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_condition;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isJump = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isJump;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isLink = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isLink;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_idx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_idx;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isIndirect = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_isIndirect;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_laCfIdx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchCtrl_laCfIdx;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_opType = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_opType;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1 = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2 = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_roundingMode = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_roundingMode;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_isIntegerDest = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_isSignedCvt = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fmaNegSrc1 = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fcmpCond = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_fpuCtrl_fcmpCond;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_csrAddr = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_csrAddr;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isWrite = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isWrite;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isRead = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isRead;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isExchange = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_isExchange;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_useUimmAsSrc = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_sysCode = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_sysCode;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_isExceptionReturn = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_isTlbOp = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_isTlbOp;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_tlbOpType = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_sysCtrl_tlbOpType;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_decodeExceptionCode;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_hasDecodeException = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_hasDecodeException;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_isMicrocode = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isMicrocode;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_microcodeEntry = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_microcodeEntry;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_isSerializing = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isSerializing;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_isBranchOrJump = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_isBranchOrJump;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_isTaken = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_isTaken;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_target = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_target;
  assign RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_wasPredicted = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_decoded_branchPrediction_wasPredicted;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_physSrc1_idx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc1_idx;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_physSrc1IsFpr = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc1IsFpr;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_physSrc2_idx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc2_idx;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_physSrc2IsFpr = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physSrc2IsFpr;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_physDest_idx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physDest_idx;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_physDestIsFpr = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_physDestIsFpr;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_oldPhysDest_idx = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_oldPhysDest_idx;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_oldPhysDestIsFpr = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_oldPhysDestIsFpr;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_allocatesPhysDest = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_allocatesPhysDest;
  assign RobAllocPlugin_logic_allocatedUops_0_rename_writesToPhysReg = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_rename_writesToPhysReg;
  assign RobAllocPlugin_logic_allocatedUops_0_uniqueId = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_uniqueId;
  assign RobAllocPlugin_logic_allocatedUops_0_dispatched = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_dispatched;
  assign RobAllocPlugin_logic_allocatedUops_0_executed = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_executed;
  assign RobAllocPlugin_logic_allocatedUops_0_hasException = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_hasException;
  assign RobAllocPlugin_logic_allocatedUops_0_exceptionCode = s2_RobAlloc_IssuePipelineSignals_RENAMED_UOPS_0_exceptionCode;
  assign RobAllocPlugin_logic_allocatedUops_0_robPtr = ROBPlugin_robComponent_io_allocate_0_robPtr;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc = RobAllocPlugin_logic_allocatedUops_0_decoded_pc;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid = RobAllocPlugin_logic_allocatedUops_0_decoded_isValid;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode = RobAllocPlugin_logic_allocatedUops_0_decoded_uopCode;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit = RobAllocPlugin_logic_allocatedUops_0_decoded_exeUnit;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa = RobAllocPlugin_logic_allocatedUops_0_decoded_isa;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx = RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_idx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype = RobAllocPlugin_logic_allocatedUops_0_decoded_archDest_rtype;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn = RobAllocPlugin_logic_allocatedUops_0_decoded_writeArchDestEn;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx = RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_idx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype = RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc1_rtype;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1 = RobAllocPlugin_logic_allocatedUops_0_decoded_useArchSrc1;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx = RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_idx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype = RobAllocPlugin_logic_allocatedUops_0_decoded_archSrc2_rtype;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2 = RobAllocPlugin_logic_allocatedUops_0_decoded_useArchSrc2;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr = RobAllocPlugin_logic_allocatedUops_0_decoded_usePcForAddr;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm = RobAllocPlugin_logic_allocatedUops_0_decoded_imm;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage = RobAllocPlugin_logic_allocatedUops_0_decoded_immUsage;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid = RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_valid;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub = RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isSub;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd = RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isAdd;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned = RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_isSigned;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp = RobAllocPlugin_logic_allocatedUops_0_decoded_aluCtrl_logicOp;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid = RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_valid;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight = RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isRight;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic = RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isArithmetic;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate = RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isRotate;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord = RobAllocPlugin_logic_allocatedUops_0_decoded_shiftCtrl_isDoubleWord;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid = RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_valid;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv = RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isDiv;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned = RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isSigned;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp = RobAllocPlugin_logic_allocatedUops_0_decoded_mulDivCtrl_isWordOp;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_size;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isSignedLoad;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isStore;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isLoadLinked;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isStoreCond;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_atomicOp;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isFence;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_fenceMode;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isCacheOp;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_cacheOpType;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch = RobAllocPlugin_logic_allocatedUops_0_decoded_memCtrl_isPrefetch;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition = RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_condition;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump = RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isJump;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink = RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isLink;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx = RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_idx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype = RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_linkReg_rtype;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect = RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_isIndirect;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx = RobAllocPlugin_logic_allocatedUops_0_decoded_branchCtrl_laCfIdx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_opType;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1 = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc1;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2 = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeSrc2;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fpSizeDest;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_roundingMode;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_isIntegerDest;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_isSignedCvt;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1 = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fmaNegSrc1;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond = RobAllocPlugin_logic_allocatedUops_0_decoded_fpuCtrl_fcmpCond;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr = RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_csrAddr;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite = RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isWrite;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead = RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isRead;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange = RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_isExchange;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc = RobAllocPlugin_logic_allocatedUops_0_decoded_csrCtrl_useUimmAsSrc;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode = RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_sysCode;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn = RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_isExceptionReturn;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp = RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_isTlbOp;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType = RobAllocPlugin_logic_allocatedUops_0_decoded_sysCtrl_tlbOpType;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode = RobAllocPlugin_logic_allocatedUops_0_decoded_decodeExceptionCode;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException = RobAllocPlugin_logic_allocatedUops_0_decoded_hasDecodeException;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode = RobAllocPlugin_logic_allocatedUops_0_decoded_isMicrocode;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry = RobAllocPlugin_logic_allocatedUops_0_decoded_microcodeEntry;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing = RobAllocPlugin_logic_allocatedUops_0_decoded_isSerializing;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump = RobAllocPlugin_logic_allocatedUops_0_decoded_isBranchOrJump;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken = RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_isTaken;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target = RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_target;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted = RobAllocPlugin_logic_allocatedUops_0_decoded_branchPrediction_wasPredicted;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx = RobAllocPlugin_logic_allocatedUops_0_rename_physSrc1_idx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr = RobAllocPlugin_logic_allocatedUops_0_rename_physSrc1IsFpr;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx = RobAllocPlugin_logic_allocatedUops_0_rename_physSrc2_idx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr = RobAllocPlugin_logic_allocatedUops_0_rename_physSrc2IsFpr;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx = RobAllocPlugin_logic_allocatedUops_0_rename_physDest_idx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr = RobAllocPlugin_logic_allocatedUops_0_rename_physDestIsFpr;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx = RobAllocPlugin_logic_allocatedUops_0_rename_oldPhysDest_idx;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr = RobAllocPlugin_logic_allocatedUops_0_rename_oldPhysDestIsFpr;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest = RobAllocPlugin_logic_allocatedUops_0_rename_allocatesPhysDest;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg = RobAllocPlugin_logic_allocatedUops_0_rename_writesToPhysReg;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr = RobAllocPlugin_logic_allocatedUops_0_robPtr;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId = RobAllocPlugin_logic_allocatedUops_0_uniqueId;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched = RobAllocPlugin_logic_allocatedUops_0_dispatched;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_executed = RobAllocPlugin_logic_allocatedUops_0_executed;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException = RobAllocPlugin_logic_allocatedUops_0_hasException;
  assign s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode = RobAllocPlugin_logic_allocatedUops_0_exceptionCode;
  assign DispatchPlugin_logic_iqRegs_0_1_ready = issueQueueComponent_4_io_allocateIn_ready;
  assign DispatchPlugin_logic_iqRegs_1_1_ready = issueQueueComponent_5_io_allocateIn_ready;
  assign DispatchPlugin_logic_iqRegs_2_1_ready = issueQueueComponent_6_io_allocateIn_ready;
  assign DispatchPlugin_logic_iqRegs_3_1_ready = issueQueueComponent_7_io_allocateIn_ready;
  assign AluIntEU_AluIntEuPlugin_euInputPort_valid = issueQueueComponent_4_io_issueOut_valid;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_robPtr = issueQueueComponent_4_io_issueOut_payload_robPtr;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_physDest_idx = issueQueueComponent_4_io_issueOut_payload_physDest_idx;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_physDestIsFpr = issueQueueComponent_4_io_issueOut_payload_physDestIsFpr;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_writesToPhysReg = issueQueueComponent_4_io_issueOut_payload_writesToPhysReg;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_useSrc1 = issueQueueComponent_4_io_issueOut_payload_useSrc1;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Data = issueQueueComponent_4_io_issueOut_payload_src1Data;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Tag = issueQueueComponent_4_io_issueOut_payload_src1Tag;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Ready = issueQueueComponent_4_io_issueOut_payload_src1Ready;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_src1IsFpr = issueQueueComponent_4_io_issueOut_payload_src1IsFpr;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_useSrc2 = issueQueueComponent_4_io_issueOut_payload_useSrc2;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Data = issueQueueComponent_4_io_issueOut_payload_src2Data;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Tag = issueQueueComponent_4_io_issueOut_payload_src2Tag;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Ready = issueQueueComponent_4_io_issueOut_payload_src2Ready;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_src2IsFpr = issueQueueComponent_4_io_issueOut_payload_src2IsFpr;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_valid = issueQueueComponent_4_io_issueOut_payload_aluCtrl_valid;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isSub = issueQueueComponent_4_io_issueOut_payload_aluCtrl_isSub;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isAdd = issueQueueComponent_4_io_issueOut_payload_aluCtrl_isAdd;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isSigned = issueQueueComponent_4_io_issueOut_payload_aluCtrl_isSigned;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp = issueQueueComponent_4_io_issueOut_payload_aluCtrl_logicOp;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_valid = issueQueueComponent_4_io_issueOut_payload_shiftCtrl_valid;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isRight = issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isRight;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isArithmetic = issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isArithmetic;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isRotate = issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isRotate;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isDoubleWord = issueQueueComponent_4_io_issueOut_payload_shiftCtrl_isDoubleWord;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_imm = issueQueueComponent_4_io_issueOut_payload_imm;
  assign AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage = issueQueueComponent_4_io_issueOut_payload_immUsage;
  assign AluIntEU_AluIntEuPlugin_euInputPort_fire = (AluIntEU_AluIntEuPlugin_euInputPort_valid && AluIntEU_AluIntEuPlugin_euInputPort_ready);
  assign MulEU_MulEuPlugin_euInputPort_valid = issueQueueComponent_5_io_issueOut_valid;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_pc = issueQueueComponent_5_io_issueOut_payload_uop_decoded_pc;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isValid = issueQueueComponent_5_io_issueOut_payload_uop_decoded_isValid;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_uopCode = issueQueueComponent_5_io_issueOut_payload_uop_decoded_uopCode;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_exeUnit = issueQueueComponent_5_io_issueOut_payload_uop_decoded_exeUnit;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isa = issueQueueComponent_5_io_issueOut_payload_uop_decoded_isa;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_idx = issueQueueComponent_5_io_issueOut_payload_uop_decoded_archDest_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archDest_rtype = issueQueueComponent_5_io_issueOut_payload_uop_decoded_archDest_rtype;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_writeArchDestEn = issueQueueComponent_5_io_issueOut_payload_uop_decoded_writeArchDestEn;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_idx = issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc1_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc1_rtype = issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc1_rtype;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_useArchSrc1 = issueQueueComponent_5_io_issueOut_payload_uop_decoded_useArchSrc1;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_idx = issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc2_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_archSrc2_rtype = issueQueueComponent_5_io_issueOut_payload_uop_decoded_archSrc2_rtype;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_useArchSrc2 = issueQueueComponent_5_io_issueOut_payload_uop_decoded_useArchSrc2;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_usePcForAddr = issueQueueComponent_5_io_issueOut_payload_uop_decoded_usePcForAddr;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_imm = issueQueueComponent_5_io_issueOut_payload_uop_decoded_imm;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_immUsage = issueQueueComponent_5_io_issueOut_payload_uop_decoded_immUsage;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_valid = issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_valid;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_isSub = issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isSub;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_isAdd = issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isAdd;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_isSigned = issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_isSigned;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_aluCtrl_logicOp = issueQueueComponent_5_io_issueOut_payload_uop_decoded_aluCtrl_logicOp;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_valid = issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_valid;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_isRight = issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isRight;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_isArithmetic = issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_isRotate = issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_shiftCtrl_isDoubleWord = issueQueueComponent_5_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_mulDivCtrl_valid = issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_valid;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_mulDivCtrl_isDiv = issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_mulDivCtrl_isSigned = issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_mulDivCtrl_isWordOp = issueQueueComponent_5_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_size = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_size;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isSignedLoad = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isStore = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isStore;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isLoadLinked = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isStoreCond = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_atomicOp = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_atomicOp;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isFence = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isFence;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_fenceMode = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_fenceMode;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isCacheOp = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_cacheOpType = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_memCtrl_isPrefetch = issueQueueComponent_5_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_condition = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_condition;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_isJump = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isJump;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_isLink = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isLink;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_idx = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_linkReg_rtype = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_isIndirect = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchCtrl_laCfIdx = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_opType = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_opType;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fpSizeDest = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_roundingMode = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_isIntegerDest = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_isSignedCvt = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_fpuCtrl_fcmpCond = issueQueueComponent_5_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_csrAddr = issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_isWrite = issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isWrite;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_isRead = issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isRead;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_isExchange = issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_isExchange;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_csrCtrl_useUimmAsSrc = issueQueueComponent_5_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_sysCtrl_sysCode = issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_sysCode;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_sysCtrl_isExceptionReturn = issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_sysCtrl_isTlbOp = issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_sysCtrl_tlbOpType = issueQueueComponent_5_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_decodeExceptionCode = issueQueueComponent_5_io_issueOut_payload_uop_decoded_decodeExceptionCode;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_hasDecodeException = issueQueueComponent_5_io_issueOut_payload_uop_decoded_hasDecodeException;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isMicrocode = issueQueueComponent_5_io_issueOut_payload_uop_decoded_isMicrocode;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_microcodeEntry = issueQueueComponent_5_io_issueOut_payload_uop_decoded_microcodeEntry;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isSerializing = issueQueueComponent_5_io_issueOut_payload_uop_decoded_isSerializing;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_isBranchOrJump = issueQueueComponent_5_io_issueOut_payload_uop_decoded_isBranchOrJump;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchPrediction_isTaken = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_isTaken;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchPrediction_target = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_target;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_decoded_branchPrediction_wasPredicted = issueQueueComponent_5_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physSrc1_idx = issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc1_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physSrc1IsFpr = issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc1IsFpr;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physSrc2_idx = issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc2_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physSrc2IsFpr = issueQueueComponent_5_io_issueOut_payload_uop_rename_physSrc2IsFpr;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physDest_idx = issueQueueComponent_5_io_issueOut_payload_uop_rename_physDest_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_physDestIsFpr = issueQueueComponent_5_io_issueOut_payload_uop_rename_physDestIsFpr;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_oldPhysDest_idx = issueQueueComponent_5_io_issueOut_payload_uop_rename_oldPhysDest_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_oldPhysDestIsFpr = issueQueueComponent_5_io_issueOut_payload_uop_rename_oldPhysDestIsFpr;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_allocatesPhysDest = issueQueueComponent_5_io_issueOut_payload_uop_rename_allocatesPhysDest;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_rename_writesToPhysReg = issueQueueComponent_5_io_issueOut_payload_uop_rename_writesToPhysReg;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_robPtr = issueQueueComponent_5_io_issueOut_payload_uop_robPtr;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_uniqueId = issueQueueComponent_5_io_issueOut_payload_uop_uniqueId;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_dispatched = issueQueueComponent_5_io_issueOut_payload_uop_dispatched;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_executed = issueQueueComponent_5_io_issueOut_payload_uop_executed;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_hasException = issueQueueComponent_5_io_issueOut_payload_uop_hasException;
  assign MulEU_MulEuPlugin_euInputPort_payload_uop_exceptionCode = issueQueueComponent_5_io_issueOut_payload_uop_exceptionCode;
  assign MulEU_MulEuPlugin_euInputPort_payload_robPtr = issueQueueComponent_5_io_issueOut_payload_robPtr;
  assign MulEU_MulEuPlugin_euInputPort_payload_physDest_idx = issueQueueComponent_5_io_issueOut_payload_physDest_idx;
  assign MulEU_MulEuPlugin_euInputPort_payload_physDestIsFpr = issueQueueComponent_5_io_issueOut_payload_physDestIsFpr;
  assign MulEU_MulEuPlugin_euInputPort_payload_writesToPhysReg = issueQueueComponent_5_io_issueOut_payload_writesToPhysReg;
  assign MulEU_MulEuPlugin_euInputPort_payload_useSrc1 = issueQueueComponent_5_io_issueOut_payload_useSrc1;
  assign MulEU_MulEuPlugin_euInputPort_payload_src1Data = issueQueueComponent_5_io_issueOut_payload_src1Data;
  assign MulEU_MulEuPlugin_euInputPort_payload_src1Tag = issueQueueComponent_5_io_issueOut_payload_src1Tag;
  assign MulEU_MulEuPlugin_euInputPort_payload_src1Ready = issueQueueComponent_5_io_issueOut_payload_src1Ready;
  assign MulEU_MulEuPlugin_euInputPort_payload_src1IsFpr = issueQueueComponent_5_io_issueOut_payload_src1IsFpr;
  assign MulEU_MulEuPlugin_euInputPort_payload_useSrc2 = issueQueueComponent_5_io_issueOut_payload_useSrc2;
  assign MulEU_MulEuPlugin_euInputPort_payload_src2Data = issueQueueComponent_5_io_issueOut_payload_src2Data;
  assign MulEU_MulEuPlugin_euInputPort_payload_src2Tag = issueQueueComponent_5_io_issueOut_payload_src2Tag;
  assign MulEU_MulEuPlugin_euInputPort_payload_src2Ready = issueQueueComponent_5_io_issueOut_payload_src2Ready;
  assign MulEU_MulEuPlugin_euInputPort_payload_src2IsFpr = issueQueueComponent_5_io_issueOut_payload_src2IsFpr;
  assign MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_valid = issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_valid;
  assign MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isDiv = issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isDiv;
  assign MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isSigned = issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isSigned;
  assign MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isWordOp = issueQueueComponent_5_io_issueOut_payload_mulDivCtrl_isWordOp;
  assign MulEU_MulEuPlugin_euInputPort_fire = (MulEU_MulEuPlugin_euInputPort_valid && MulEU_MulEuPlugin_euInputPort_ready);
  assign BranchEU_BranchEuPlugin_euInputPort_valid = issueQueueComponent_6_io_issueOut_valid;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_robPtr = issueQueueComponent_6_io_issueOut_payload_robPtr;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_physDest_idx = issueQueueComponent_6_io_issueOut_payload_physDest_idx;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_physDestIsFpr = issueQueueComponent_6_io_issueOut_payload_physDestIsFpr;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_writesToPhysReg = issueQueueComponent_6_io_issueOut_payload_writesToPhysReg;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_useSrc1 = issueQueueComponent_6_io_issueOut_payload_useSrc1;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_src1Data = issueQueueComponent_6_io_issueOut_payload_src1Data;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_src1Tag = issueQueueComponent_6_io_issueOut_payload_src1Tag;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_src1Ready = issueQueueComponent_6_io_issueOut_payload_src1Ready;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_src1IsFpr = issueQueueComponent_6_io_issueOut_payload_src1IsFpr;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_useSrc2 = issueQueueComponent_6_io_issueOut_payload_useSrc2;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_src2Data = issueQueueComponent_6_io_issueOut_payload_src2Data;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_src2Tag = issueQueueComponent_6_io_issueOut_payload_src2Tag;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_src2Ready = issueQueueComponent_6_io_issueOut_payload_src2Ready;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_src2IsFpr = issueQueueComponent_6_io_issueOut_payload_src2IsFpr;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition = issueQueueComponent_6_io_issueOut_payload_branchCtrl_condition;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isJump = issueQueueComponent_6_io_issueOut_payload_branchCtrl_isJump;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isLink = issueQueueComponent_6_io_issueOut_payload_branchCtrl_isLink;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_idx = issueQueueComponent_6_io_issueOut_payload_branchCtrl_linkReg_idx;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype = issueQueueComponent_6_io_issueOut_payload_branchCtrl_linkReg_rtype;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isIndirect = issueQueueComponent_6_io_issueOut_payload_branchCtrl_isIndirect;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_laCfIdx = issueQueueComponent_6_io_issueOut_payload_branchCtrl_laCfIdx;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_imm = issueQueueComponent_6_io_issueOut_payload_imm;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_pc = issueQueueComponent_6_io_issueOut_payload_pc;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_isTaken = issueQueueComponent_6_io_issueOut_payload_branchPrediction_isTaken;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_target = issueQueueComponent_6_io_issueOut_payload_branchPrediction_target;
  assign BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_wasPredicted = issueQueueComponent_6_io_issueOut_payload_branchPrediction_wasPredicted;
  assign BranchEU_BranchEuPlugin_euInputPort_fire = (BranchEU_BranchEuPlugin_euInputPort_valid && BranchEU_BranchEuPlugin_euInputPort_ready);
  assign LsuEU_LsuEuPlugin_euInputPort_valid = issueQueueComponent_7_io_issueOut_valid;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_robPtr = issueQueueComponent_7_io_issueOut_payload_robPtr;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_physDest_idx = issueQueueComponent_7_io_issueOut_payload_physDest_idx;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_physDestIsFpr = issueQueueComponent_7_io_issueOut_payload_physDestIsFpr;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_writesToPhysReg = issueQueueComponent_7_io_issueOut_payload_writesToPhysReg;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_useSrc1 = issueQueueComponent_7_io_issueOut_payload_useSrc1;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_src1Data = issueQueueComponent_7_io_issueOut_payload_src1Data;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_src1Tag = issueQueueComponent_7_io_issueOut_payload_src1Tag;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_src1Ready = issueQueueComponent_7_io_issueOut_payload_src1Ready;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_src1IsFpr = issueQueueComponent_7_io_issueOut_payload_src1IsFpr;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_useSrc2 = issueQueueComponent_7_io_issueOut_payload_useSrc2;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_src2Data = issueQueueComponent_7_io_issueOut_payload_src2Data;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_src2Tag = issueQueueComponent_7_io_issueOut_payload_src2Tag;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_src2Ready = issueQueueComponent_7_io_issueOut_payload_src2Ready;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_src2IsFpr = issueQueueComponent_7_io_issueOut_payload_src2IsFpr;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size = issueQueueComponent_7_io_issueOut_payload_memCtrl_size;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isSignedLoad = issueQueueComponent_7_io_issueOut_payload_memCtrl_isSignedLoad;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isStore = issueQueueComponent_7_io_issueOut_payload_memCtrl_isStore;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isLoadLinked = issueQueueComponent_7_io_issueOut_payload_memCtrl_isLoadLinked;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isStoreCond = issueQueueComponent_7_io_issueOut_payload_memCtrl_isStoreCond;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_atomicOp = issueQueueComponent_7_io_issueOut_payload_memCtrl_atomicOp;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isFence = issueQueueComponent_7_io_issueOut_payload_memCtrl_isFence;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_fenceMode = issueQueueComponent_7_io_issueOut_payload_memCtrl_fenceMode;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isCacheOp = issueQueueComponent_7_io_issueOut_payload_memCtrl_isCacheOp;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_cacheOpType = issueQueueComponent_7_io_issueOut_payload_memCtrl_cacheOpType;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isPrefetch = issueQueueComponent_7_io_issueOut_payload_memCtrl_isPrefetch;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_imm = issueQueueComponent_7_io_issueOut_payload_imm;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_usePc = issueQueueComponent_7_io_issueOut_payload_usePc;
  assign LsuEU_LsuEuPlugin_euInputPort_payload_pcData = issueQueueComponent_7_io_issueOut_payload_pcData;
  assign LsuEU_LsuEuPlugin_euInputPort_fire = (LsuEU_LsuEuPlugin_euInputPort_valid && LsuEU_LsuEuPlugin_euInputPort_ready);
  assign oneShot_20_io_triggerIn = (AluIntEU_AluIntEuPlugin_euInputPort_fire && (_zz_when_Debug_l71 < _zz_io_triggerIn_12));
  assign _zz_when_Debug_l71_7 = 5'h17;
  assign when_Debug_l71_6 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_6_1);
  assign DispatchPlugin_logic_physSrc1ConflictS1 = 1'b0;
  assign DispatchPlugin_logic_physSrc1ConflictS2 = ((s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid && s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest) && (s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx == s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx));
  assign DispatchPlugin_logic_physSrc2ConflictS1 = 1'b0;
  assign DispatchPlugin_logic_physSrc2ConflictS2 = ((s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid && s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest) && (s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx == s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx));
  assign DispatchPlugin_logic_src1SetBypass = (DispatchPlugin_logic_physSrc1ConflictS1 || DispatchPlugin_logic_physSrc1ConflictS2);
  assign DispatchPlugin_logic_src2SetBypass = (DispatchPlugin_logic_physSrc2ConflictS1 || DispatchPlugin_logic_physSrc2ConflictS2);
  assign DispatchPlugin_logic_src1ReadyCandidate = ((! BusyTablePlugin_early_setup_busyTableReg[s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx]) || BusyTablePlugin_early_setup_clearMask[s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx]);
  assign DispatchPlugin_logic_src1InitialReady = ((! s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1) || (DispatchPlugin_logic_src1ReadyCandidate && (! DispatchPlugin_logic_src1SetBypass)));
  assign DispatchPlugin_logic_src2ReadyCandidate = ((! BusyTablePlugin_early_setup_busyTableReg[s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx]) || BusyTablePlugin_early_setup_clearMask[s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx]);
  assign DispatchPlugin_logic_src2InitialReady = ((! s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2) || (DispatchPlugin_logic_src2ReadyCandidate && (! DispatchPlugin_logic_src2SetBypass)));
  assign DispatchPlugin_logic_dispatchOH = {(|{(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_3_0_1),(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_3_0_0)}),{(|{(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_2_0_2),{_zz_DispatchPlugin_logic_dispatchOH,_zz_DispatchPlugin_logic_dispatchOH_1}}),{(|(s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode == DispatchPlugin_logic_iqRegs_1_0_0)),(|{_zz_DispatchPlugin_logic_dispatchOH_2,{_zz_DispatchPlugin_logic_dispatchOH_3,_zz_DispatchPlugin_logic_dispatchOH_4}})}}};
  assign _zz_DispatchPlugin_logic_destinationIqReady = DispatchPlugin_logic_dispatchOH[3];
  assign _zz_DispatchPlugin_logic_destinationIqReady_1 = (DispatchPlugin_logic_dispatchOH[1] || _zz_DispatchPlugin_logic_destinationIqReady);
  assign _zz_DispatchPlugin_logic_destinationIqReady_2 = (DispatchPlugin_logic_dispatchOH[2] || _zz_DispatchPlugin_logic_destinationIqReady);
  assign DispatchPlugin_logic_destinationIqReady = _zz_DispatchPlugin_logic_destinationIqReady_3;
  assign s3_Dispatch_haltRequest_DispatchPlugin_l78 = ((s3_Dispatch_valid && s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid) && (! DispatchPlugin_logic_destinationIqReady));
  assign DispatchPlugin_logic_iqRegs_0_1_valid = ((s3_Dispatch_isFiring && s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid) && DispatchPlugin_logic_dispatchOH[0]);
  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_pc = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isValid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isValid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_uopCode = (5'bxxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_exeUnit = (4'bxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isa = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archDest_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_writeArchDestEn = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_writeArchDestEn = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc1_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_useArchSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_useArchSrc1 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_archSrc2_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_useArchSrc2 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_useArchSrc2 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_usePcForAddr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_usePcForAddr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_imm = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_imm = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_immUsage = (3'bxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isSub = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isSub = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isAdd = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isAdd = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isSigned = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_isSigned = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_aluCtrl_logicOp = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isRight = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isRight = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isArithmetic = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isArithmetic = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isRotate = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isRotate = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isDoubleWord = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_shiftCtrl_isDoubleWord = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isDiv = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isDiv = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isSigned = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isSigned = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isWordOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_mulDivCtrl_isWordOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_size = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isSignedLoad = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isSignedLoad = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isStore = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isStore = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isLoadLinked = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isLoadLinked = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isStoreCond = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isStoreCond = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_atomicOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_atomicOp = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isFence = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isFence = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_fenceMode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_fenceMode = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isCacheOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isCacheOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_cacheOpType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_cacheOpType = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isPrefetch = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_memCtrl_isPrefetch = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_condition = (5'bxxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isJump = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isJump = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isLink = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isLink = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_linkReg_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isIndirect = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_isIndirect = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_laCfIdx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchCtrl_laCfIdx = 3'bxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_opType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_opType = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fpSizeDest = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_roundingMode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_roundingMode = 3'bxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_isIntegerDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_isIntegerDest = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_isSignedCvt = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_isSignedCvt = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fcmpCond = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_fpuCtrl_fcmpCond = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_csrAddr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_csrAddr = 14'bxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isWrite = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isWrite = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isRead = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isRead = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isExchange = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_isExchange = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_useUimmAsSrc = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_csrCtrl_useUimmAsSrc = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_sysCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_sysCode = 20'bxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_isExceptionReturn = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_isExceptionReturn = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_isTlbOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_isTlbOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_tlbOpType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_sysCtrl_tlbOpType = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_decodeExceptionCode = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_hasDecodeException = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_hasDecodeException = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isMicrocode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isMicrocode = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_microcodeEntry = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_microcodeEntry = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isSerializing = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isSerializing = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isBranchOrJump = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_isBranchOrJump = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_isTaken = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_isTaken = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_target = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_wasPredicted = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_decoded_branchPrediction_wasPredicted = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc1_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc1_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc1IsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc1IsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc2_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc2_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc2IsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physSrc2IsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physDest_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physDestIsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_physDestIsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_oldPhysDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_oldPhysDest_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_oldPhysDestIsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_oldPhysDestIsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_allocatesPhysDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_allocatesPhysDest = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_writesToPhysReg = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_rename_writesToPhysReg = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_robPtr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_robPtr = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_uniqueId = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_uniqueId = 16'bxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_dispatched = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_dispatched = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_executed = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_executed;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_executed = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_hasException = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_hasException = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_exceptionCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_uop_exceptionCode = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_src1InitialReady = DispatchPlugin_logic_src1InitialReady;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_src1InitialReady = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_0_1_valid) begin
      DispatchPlugin_logic_iqRegs_0_1_payload_src2InitialReady = DispatchPlugin_logic_src2InitialReady;
    end else begin
      DispatchPlugin_logic_iqRegs_0_1_payload_src2InitialReady = 1'bx;
    end
  end

  assign DispatchPlugin_logic_iqRegs_1_1_valid = ((s3_Dispatch_isFiring && s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid) && DispatchPlugin_logic_dispatchOH[1]);
  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_pc = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isValid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isValid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_uopCode = (5'bxxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_exeUnit = (4'bxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isa = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archDest_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_writeArchDestEn = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_writeArchDestEn = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc1_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_useArchSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_useArchSrc1 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_archSrc2_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_useArchSrc2 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_useArchSrc2 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_usePcForAddr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_usePcForAddr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_imm = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_imm = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_immUsage = (3'bxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isSub = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isSub = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isAdd = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isAdd = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isSigned = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_isSigned = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_aluCtrl_logicOp = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isRight = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isRight = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isArithmetic = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isArithmetic = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isRotate = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isRotate = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isDoubleWord = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_shiftCtrl_isDoubleWord = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isDiv = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isDiv = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isSigned = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isSigned = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isWordOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_mulDivCtrl_isWordOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_size = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isSignedLoad = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isSignedLoad = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isStore = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isStore = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isLoadLinked = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isLoadLinked = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isStoreCond = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isStoreCond = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_atomicOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_atomicOp = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isFence = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isFence = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_fenceMode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_fenceMode = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isCacheOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isCacheOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_cacheOpType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_cacheOpType = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isPrefetch = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_memCtrl_isPrefetch = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_condition = (5'bxxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isJump = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isJump = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isLink = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isLink = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_linkReg_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isIndirect = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_isIndirect = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_laCfIdx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchCtrl_laCfIdx = 3'bxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_opType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_opType = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fpSizeDest = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_roundingMode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_roundingMode = 3'bxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_isIntegerDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_isIntegerDest = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_isSignedCvt = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_isSignedCvt = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fcmpCond = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_fpuCtrl_fcmpCond = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_csrAddr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_csrAddr = 14'bxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isWrite = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isWrite = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isRead = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isRead = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isExchange = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_isExchange = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_useUimmAsSrc = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_csrCtrl_useUimmAsSrc = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_sysCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_sysCode = 20'bxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_isExceptionReturn = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_isExceptionReturn = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_isTlbOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_isTlbOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_tlbOpType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_sysCtrl_tlbOpType = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_decodeExceptionCode = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_hasDecodeException = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_hasDecodeException = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isMicrocode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isMicrocode = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_microcodeEntry = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_microcodeEntry = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isSerializing = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isSerializing = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isBranchOrJump = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_isBranchOrJump = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_isTaken = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_isTaken = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_target = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_wasPredicted = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_decoded_branchPrediction_wasPredicted = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc1_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc1_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc1IsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc1IsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc2_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc2_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc2IsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physSrc2IsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physDest_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physDestIsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_physDestIsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_oldPhysDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_oldPhysDest_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_oldPhysDestIsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_oldPhysDestIsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_allocatesPhysDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_allocatesPhysDest = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_writesToPhysReg = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_rename_writesToPhysReg = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_robPtr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_robPtr = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_uniqueId = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_uniqueId = 16'bxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_dispatched = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_dispatched = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_executed = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_executed;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_executed = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_hasException = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_hasException = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_exceptionCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_uop_exceptionCode = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_src1InitialReady = DispatchPlugin_logic_src1InitialReady;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_src1InitialReady = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_1_1_valid) begin
      DispatchPlugin_logic_iqRegs_1_1_payload_src2InitialReady = DispatchPlugin_logic_src2InitialReady;
    end else begin
      DispatchPlugin_logic_iqRegs_1_1_payload_src2InitialReady = 1'bx;
    end
  end

  assign DispatchPlugin_logic_iqRegs_2_1_valid = ((s3_Dispatch_isFiring && s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid) && DispatchPlugin_logic_dispatchOH[2]);
  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_pc = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isValid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isValid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_uopCode = (5'bxxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_exeUnit = (4'bxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isa = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archDest_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_writeArchDestEn = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_writeArchDestEn = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc1_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_useArchSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_useArchSrc1 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_archSrc2_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_useArchSrc2 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_useArchSrc2 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_usePcForAddr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_usePcForAddr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_imm = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_imm = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_immUsage = (3'bxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isSub = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isSub = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isAdd = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isAdd = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isSigned = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_isSigned = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_aluCtrl_logicOp = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isRight = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isRight = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isArithmetic = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isArithmetic = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isRotate = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isRotate = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isDoubleWord = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_shiftCtrl_isDoubleWord = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isDiv = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isDiv = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isSigned = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isSigned = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isWordOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_mulDivCtrl_isWordOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_size = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isSignedLoad = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isSignedLoad = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isStore = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isStore = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isLoadLinked = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isLoadLinked = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isStoreCond = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isStoreCond = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_atomicOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_atomicOp = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isFence = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isFence = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_fenceMode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_fenceMode = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isCacheOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isCacheOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_cacheOpType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_cacheOpType = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isPrefetch = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_memCtrl_isPrefetch = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_condition = (5'bxxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isJump = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isJump = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isLink = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isLink = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_linkReg_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isIndirect = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_isIndirect = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_laCfIdx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchCtrl_laCfIdx = 3'bxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_opType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_opType = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fpSizeDest = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_roundingMode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_roundingMode = 3'bxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_isIntegerDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_isIntegerDest = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_isSignedCvt = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_isSignedCvt = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fcmpCond = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_fpuCtrl_fcmpCond = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_csrAddr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_csrAddr = 14'bxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isWrite = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isWrite = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isRead = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isRead = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isExchange = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_isExchange = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_useUimmAsSrc = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_csrCtrl_useUimmAsSrc = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_sysCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_sysCode = 20'bxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_isExceptionReturn = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_isExceptionReturn = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_isTlbOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_isTlbOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_tlbOpType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_sysCtrl_tlbOpType = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_decodeExceptionCode = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_hasDecodeException = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_hasDecodeException = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isMicrocode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isMicrocode = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_microcodeEntry = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_microcodeEntry = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isSerializing = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isSerializing = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isBranchOrJump = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_isBranchOrJump = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_isTaken = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_isTaken = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_target = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_wasPredicted = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_decoded_branchPrediction_wasPredicted = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc1_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc1_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc1IsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc1IsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc2_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc2_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc2IsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physSrc2IsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physDest_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physDestIsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_physDestIsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_oldPhysDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_oldPhysDest_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_oldPhysDestIsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_oldPhysDestIsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_allocatesPhysDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_allocatesPhysDest = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_writesToPhysReg = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_rename_writesToPhysReg = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_robPtr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_robPtr = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_uniqueId = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_uniqueId = 16'bxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_dispatched = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_dispatched = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_executed = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_executed;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_executed = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_hasException = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_hasException = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_exceptionCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_uop_exceptionCode = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_src1InitialReady = DispatchPlugin_logic_src1InitialReady;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_src1InitialReady = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_2_1_valid) begin
      DispatchPlugin_logic_iqRegs_2_1_payload_src2InitialReady = DispatchPlugin_logic_src2InitialReady;
    end else begin
      DispatchPlugin_logic_iqRegs_2_1_payload_src2InitialReady = 1'bx;
    end
  end

  assign DispatchPlugin_logic_iqRegs_3_1_valid = ((s3_Dispatch_isFiring && s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid) && DispatchPlugin_logic_dispatchOH[3]);
  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_pc = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isValid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isValid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_uopCode = (5'bxxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_exeUnit = (4'bxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isa = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archDest_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_writeArchDestEn = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_writeArchDestEn = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc1_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_useArchSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_useArchSrc1 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_archSrc2_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_useArchSrc2 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_useArchSrc2 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_usePcForAddr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_usePcForAddr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_imm = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_imm = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_immUsage = (3'bxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isSub = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isSub = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isAdd = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isAdd = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isSigned = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_isSigned = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_aluCtrl_logicOp = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isRight = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isRight = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isArithmetic = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isArithmetic = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isRotate = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isRotate = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isDoubleWord = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_shiftCtrl_isDoubleWord = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_valid = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_valid = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isDiv = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isDiv = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isSigned = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isSigned = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isWordOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_mulDivCtrl_isWordOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_size = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isSignedLoad = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isSignedLoad = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isStore = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isStore = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isLoadLinked = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isLoadLinked = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isStoreCond = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isStoreCond = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_atomicOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_atomicOp = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isFence = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isFence = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_fenceMode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_fenceMode = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isCacheOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isCacheOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_cacheOpType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_cacheOpType = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isPrefetch = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_memCtrl_isPrefetch = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_condition = (5'bxxxxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isJump = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isJump = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isLink = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isLink = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_idx = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_linkReg_rtype = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isIndirect = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_isIndirect = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_laCfIdx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchCtrl_laCfIdx = 3'bxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_opType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_opType = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fpSizeDest = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_roundingMode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_roundingMode = 3'bxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_isIntegerDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_isIntegerDest = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_isSignedCvt = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_isSignedCvt = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fcmpCond = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_fpuCtrl_fcmpCond = 5'bxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_csrAddr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_csrAddr = 14'bxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isWrite = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isWrite = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isRead = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isRead = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isExchange = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_isExchange = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_useUimmAsSrc = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_csrCtrl_useUimmAsSrc = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_sysCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_sysCode = 20'bxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_isExceptionReturn = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_isExceptionReturn = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_isTlbOp = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_isTlbOp = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_tlbOpType = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_sysCtrl_tlbOpType = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_decodeExceptionCode = (2'bxx);
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_hasDecodeException = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_hasDecodeException = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isMicrocode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isMicrocode = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_microcodeEntry = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_microcodeEntry = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isSerializing = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isSerializing = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isBranchOrJump = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_isBranchOrJump = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_isTaken = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_isTaken = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_target = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_wasPredicted = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_decoded_branchPrediction_wasPredicted = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc1_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc1_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc1IsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc1IsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc2_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc2_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc2IsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physSrc2IsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physDest_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physDestIsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_physDestIsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_oldPhysDest_idx = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_oldPhysDest_idx = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_oldPhysDestIsFpr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_oldPhysDestIsFpr = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_allocatesPhysDest = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_allocatesPhysDest = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_writesToPhysReg = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_rename_writesToPhysReg = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_robPtr = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_robPtr = 4'bxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_uniqueId = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_uniqueId = 16'bxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_dispatched = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_dispatched = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_executed = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_executed;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_executed = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_hasException = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_hasException = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_exceptionCode = s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_uop_exceptionCode = 8'bxxxxxxxx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_src1InitialReady = DispatchPlugin_logic_src1InitialReady;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_src1InitialReady = 1'bx;
    end
  end

  always @(*) begin
    if(DispatchPlugin_logic_iqRegs_3_1_valid) begin
      DispatchPlugin_logic_iqRegs_3_1_payload_src2InitialReady = DispatchPlugin_logic_src2InitialReady;
    end else begin
      DispatchPlugin_logic_iqRegs_3_1_payload_src2InitialReady = 1'bx;
    end
  end

  assign when_DispatchPlugin_l100 = (s3_Dispatch_isFiring && s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid);
  assign CommitPlugin_commitEnableExt = 1'b1;
  assign CoreNSCSCCSetupPlugin_logic_instructionVec_0 = FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_instruction;
  assign CoreNSCSCCSetupPlugin_logic_instructionVec_1 = 32'h0;
  assign CoreNSCSCCSetupPlugin_logic_instructionVec_2 = 32'h0;
  assign CoreNSCSCCSetupPlugin_logic_instructionVec_3 = 32'h0;
  assign s0_Decode_valid = FetchPipelinePlugin_setup_fetchOutput_io_pop_valid;
  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_GROUP_PC_IN = FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_pc;
    end else begin
      s0_Decode_IssuePipelineSignals_GROUP_PC_IN = 32'h0;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_0 = CoreNSCSCCSetupPlugin_logic_instructionVec_0;
    end else begin
      s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_1 = CoreNSCSCCSetupPlugin_logic_instructionVec_1;
    end else begin
      s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_2 = CoreNSCSCCSetupPlugin_logic_instructionVec_2;
    end else begin
      s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_2 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_3 = CoreNSCSCCSetupPlugin_logic_instructionVec_3;
    end else begin
      s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_3 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_isTaken = FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_isTaken;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_isTaken = 1'bx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_target = FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_target;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_wasPredicted = FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_bpuPrediction_wasPredicted;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_0_wasPredicted = 1'bx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_isTaken = 1'bx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_isTaken = 1'bx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_wasPredicted = 1'bx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_1_wasPredicted = 1'bx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_isTaken = 1'bx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_isTaken = 1'bx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_wasPredicted = 1'bx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_2_wasPredicted = 1'bx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_isTaken = 1'bx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_isTaken = 1'bx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_wasPredicted = 1'bx;
    end else begin
      s0_Decode_IssuePipelineSignals_BRANCH_PREDICTION_3_wasPredicted = 1'bx;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_VALID_MASK = 4'b0001;
    end else begin
      s0_Decode_IssuePipelineSignals_VALID_MASK = 4'b0000;
    end
  end

  always @(*) begin
    if(FetchPipelinePlugin_setup_fetchOutput_io_pop_valid) begin
      s0_Decode_IssuePipelineSignals_IS_FAULT_IN = 1'b0;
    end else begin
      s0_Decode_IssuePipelineSignals_IS_FAULT_IN = 1'b0;
    end
  end

  assign DebugDisplayPlugin_hw_dpyController_io_dp0 = (! DebugDisplayPlugin_logic_displayArea_dpToggle);
  assign s0_Dispatch_valid = AluIntEU_AluIntEuPlugin_euInputPort_valid;
  assign AluIntEU_AluIntEuPlugin_euInputPort_ready = s0_Dispatch_ready_1;
  assign _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2 = AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_logicOp;
  assign _zz_io_iqEntryIn_payload_immUsage_2 = AluIntEU_AluIntEuPlugin_euInputPort_payload_immUsage;
  assign s1_ReadRegs_isFiring = (s1_ReadRegs_valid && s1_ReadRegs_ready);
  assign AluIntEU_AluIntEuPlugin_gprReadPorts_0_valid = (s1_ReadRegs_isFiring && _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_valid);
  assign AluIntEU_AluIntEuPlugin_gprReadPorts_0_address = _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_address;
  assign AluIntEU_AluIntEuPlugin_gprReadPorts_1_valid = (s1_ReadRegs_isFiring && _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_valid);
  assign AluIntEU_AluIntEuPlugin_gprReadPorts_1_address = _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_address;
  assign _zz_io_iqEntryIn_payload_src2Data_1 = ((_zz_io_iqEntryIn_payload_immUsage == ImmUsageType_SRC_ALU) ? _zz_io_iqEntryIn_payload_imm : _zz_io_iqEntryIn_payload_src2Data);
  assign _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_1 = AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_exceptionCode;
  assign s2_Execute_isFiring = (s2_Execute_valid && s2_Execute_ready);
  assign _zz_51 = _zz_io_iqEntryIn_payload_immUsage;
  assign s3_Writeback_isFiring = (s3_Writeback_valid && s3_Writeback_ready);
  assign s3_Writeback_isFlushed = ROBPlugin_aggregatedFlushSignal_valid;
  assign when_Connection_l66_1 = (|{ROBPlugin_aggregatedFlushSignal_valid,ROBPlugin_aggregatedFlushSignal_valid});
  assign s2_Execute_isFlushed = when_Connection_l66_1;
  assign when_Connection_l66_2 = (|{when_Connection_l66_1,ROBPlugin_aggregatedFlushSignal_valid});
  assign s1_ReadRegs_isFlushed = when_Connection_l66_2;
  assign s0_Dispatch_isFlushed_1 = (|{when_Connection_l66_2,ROBPlugin_aggregatedFlushSignal_valid});
  assign s0_Dispatch_isFlushingRoot_1 = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign s1_ReadRegs_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign s2_Execute_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign s3_Writeback_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  always @(*) begin
    _zz_s1_ReadRegs_valid = s0_Dispatch_valid;
    if(s0_Dispatch_isFlushingRoot_1) begin
      _zz_s1_ReadRegs_valid = 1'b0;
    end
  end

  assign s0_Dispatch_ready_1 = 1'b1;
  always @(*) begin
    _zz_s2_Execute_valid = s1_ReadRegs_valid;
    if(s1_ReadRegs_isFlushingRoot) begin
      _zz_s2_Execute_valid = 1'b0;
    end
  end

  assign s1_ReadRegs_ready = 1'b1;
  always @(*) begin
    _zz_s3_Writeback_valid = s2_Execute_valid;
    if(s2_Execute_isFlushingRoot) begin
      _zz_s3_Writeback_valid = 1'b0;
    end
  end

  assign s2_Execute_ready = 1'b1;
  assign s3_Writeback_ready = 1'b1;
  assign when_EuBasePlugin_l230 = (ROBPlugin_aggregatedFlushSignal_valid && AluIntEU_AluIntEuPlugin_euResult_valid);
  assign AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes = (AluIntEU_AluIntEuPlugin_euResult_valid && (! ROBPlugin_aggregatedFlushSignal_valid));
  assign AluIntEU_AluIntEuPlugin_logicPhase_completesSuccessfully = (AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes && (! AluIntEU_AluIntEuPlugin_euResult_hasException));
  assign oneShot_21_io_triggerIn = (AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes && (_zz_when_Debug_l71 < _zz_io_triggerIn_14));
  assign _zz_when_Debug_l71_8 = 5'h18;
  assign when_Debug_l71_7 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_7_1);
  assign AluIntEU_AluIntEuPlugin_gprWritePort_valid = ((AluIntEU_AluIntEuPlugin_logicPhase_completesSuccessfully && AluIntEU_AluIntEuPlugin_euResult_writesToPreg) && (! AluIntEU_AluIntEuPlugin_euResult_destIsFpr));
  assign AluIntEU_AluIntEuPlugin_gprWritePort_address = AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx;
  assign AluIntEU_AluIntEuPlugin_gprWritePort_data = AluIntEU_AluIntEuPlugin_euResult_data;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_valid = AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_physRegIdx = AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_physRegData = AluIntEU_AluIntEuPlugin_euResult_data;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_robPtr = AluIntEU_AluIntEuPlugin_euResult_uop_robPtr;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_isFPR = AluIntEU_AluIntEuPlugin_euResult_destIsFpr;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_hasException = AluIntEU_AluIntEuPlugin_euResult_hasException;
  assign AluIntEU_AluIntEuPlugin_bypassOutputPort_payload_exceptionCode = AluIntEU_AluIntEuPlugin_euResult_exceptionCode;
  assign AluIntEU_AluIntEuPlugin_wakeupSourcePort_valid = (AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes && AluIntEU_AluIntEuPlugin_euResult_writesToPreg);
  assign AluIntEU_AluIntEuPlugin_wakeupSourcePort_payload_physRegIdx = AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx;
  assign AluIntEU_AluIntEuPlugin_setup_clearBusyPort_valid = (AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes && AluIntEU_AluIntEuPlugin_euResult_writesToPreg);
  assign AluIntEU_AluIntEuPlugin_setup_clearBusyPort_payload = AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx;
  assign when_EuBasePlugin_l300 = ((AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes && AluIntEU_AluIntEuPlugin_euResult_writesToPreg) && (AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx < 6'h06));
  assign mul_s0_Dispatch_valid = MulEU_MulEuPlugin_euInputPort_valid;
  assign MulEU_MulEuPlugin_euInputPort_ready = mul_s0_Dispatch_ready;
  assign mul_s1_ReadRegs_isFiring = (mul_s1_ReadRegs_valid && mul_s1_ReadRegs_ready);
  assign MulEU_MulEuPlugin_gprReadPorts_0_valid = (mul_s1_ReadRegs_isFiring && _zz_MulEU_MulEuPlugin_gprReadPorts_0_valid);
  assign MulEU_MulEuPlugin_gprReadPorts_0_address = _zz_MulEU_MulEuPlugin_gprReadPorts_0_address;
  assign MulEU_MulEuPlugin_gprReadPorts_1_valid = (mul_s1_ReadRegs_isFiring && _zz_MulEU_MulEuPlugin_gprReadPorts_1_valid);
  assign MulEU_MulEuPlugin_gprReadPorts_1_address = _zz_MulEU_MulEuPlugin_gprReadPorts_1_address;
  assign _zz_A = MulEU_MulEuPlugin_gprReadPorts_0_rsp;
  assign _zz_B = MulEU_MulEuPlugin_gprReadPorts_1_rsp;
  assign multiplierBlackbox_A = _zz_A;
  assign multiplierBlackbox_B = _zz_B;
  assign _zz_MulEU_MulEuPlugin_euResult_data = multiplierBlackbox_P;
  assign mul_s2_Execute_isFiring = (mul_s2_Execute_valid && mul_s2_Execute_ready);
  assign mul_s7_Writeback_isFiring = (mul_s7_Writeback_valid && mul_s7_Writeback_ready);
  assign mul_s7_Writeback_isFlushed = ROBPlugin_aggregatedFlushSignal_valid;
  assign when_Connection_l66_3 = (|{ROBPlugin_aggregatedFlushSignal_valid,ROBPlugin_aggregatedFlushSignal_valid});
  assign mul_s6_Execute_isFlushed = when_Connection_l66_3;
  assign when_Connection_l66_4 = (|{when_Connection_l66_3,ROBPlugin_aggregatedFlushSignal_valid});
  assign mul_s5_Execute_isFlushed = when_Connection_l66_4;
  assign when_Connection_l66_5 = (|{when_Connection_l66_4,ROBPlugin_aggregatedFlushSignal_valid});
  assign mul_s4_Execute_isFlushed = when_Connection_l66_5;
  assign when_Connection_l66_6 = (|{when_Connection_l66_5,ROBPlugin_aggregatedFlushSignal_valid});
  assign mul_s3_Execute_isFlushed = when_Connection_l66_6;
  assign when_Connection_l66_7 = (|{when_Connection_l66_6,ROBPlugin_aggregatedFlushSignal_valid});
  assign mul_s2_Execute_isFlushed = when_Connection_l66_7;
  assign when_Connection_l66_8 = (|{when_Connection_l66_7,ROBPlugin_aggregatedFlushSignal_valid});
  assign mul_s1_ReadRegs_isFlushed = when_Connection_l66_8;
  assign mul_s0_Dispatch_isFlushed = (|{when_Connection_l66_8,ROBPlugin_aggregatedFlushSignal_valid});
  assign mul_s0_Dispatch_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign mul_s1_ReadRegs_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign mul_s2_Execute_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign mul_s3_Execute_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign mul_s4_Execute_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign mul_s5_Execute_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign mul_s6_Execute_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign mul_s7_Writeback_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  always @(*) begin
    _zz_mul_s1_ReadRegs_valid = mul_s0_Dispatch_valid;
    if(mul_s0_Dispatch_isFlushingRoot) begin
      _zz_mul_s1_ReadRegs_valid = 1'b0;
    end
  end

  assign mul_s0_Dispatch_ready = 1'b1;
  always @(*) begin
    _zz_mul_s2_Execute_valid = mul_s1_ReadRegs_valid;
    if(mul_s1_ReadRegs_isFlushingRoot) begin
      _zz_mul_s2_Execute_valid = 1'b0;
    end
  end

  assign mul_s1_ReadRegs_ready = 1'b1;
  always @(*) begin
    _zz_mul_s3_Execute_valid = mul_s2_Execute_valid;
    if(mul_s2_Execute_isFlushingRoot) begin
      _zz_mul_s3_Execute_valid = 1'b0;
    end
  end

  assign mul_s2_Execute_ready = 1'b1;
  always @(*) begin
    _zz_mul_s4_Execute_valid = mul_s3_Execute_valid;
    if(mul_s3_Execute_isFlushingRoot) begin
      _zz_mul_s4_Execute_valid = 1'b0;
    end
  end

  always @(*) begin
    _zz_mul_s5_Execute_valid = mul_s4_Execute_valid;
    if(mul_s4_Execute_isFlushingRoot) begin
      _zz_mul_s5_Execute_valid = 1'b0;
    end
  end

  always @(*) begin
    _zz_mul_s6_Execute_valid = mul_s5_Execute_valid;
    if(mul_s5_Execute_isFlushingRoot) begin
      _zz_mul_s6_Execute_valid = 1'b0;
    end
  end

  always @(*) begin
    _zz_mul_s7_Writeback_valid = mul_s6_Execute_valid;
    if(mul_s6_Execute_isFlushingRoot) begin
      _zz_mul_s7_Writeback_valid = 1'b0;
    end
  end

  assign mul_s7_Writeback_ready = 1'b1;
  assign when_EuBasePlugin_l230_1 = (ROBPlugin_aggregatedFlushSignal_valid && MulEU_MulEuPlugin_euResult_valid);
  assign MulEU_MulEuPlugin_logicPhase_executionCompletes = (MulEU_MulEuPlugin_euResult_valid && (! ROBPlugin_aggregatedFlushSignal_valid));
  assign MulEU_MulEuPlugin_logicPhase_completesSuccessfully = (MulEU_MulEuPlugin_logicPhase_executionCompletes && (! MulEU_MulEuPlugin_euResult_hasException));
  assign oneShot_22_io_triggerIn = (MulEU_MulEuPlugin_logicPhase_executionCompletes && (_zz_when_Debug_l71 < _zz_io_triggerIn_16));
  assign _zz_when_Debug_l71_9 = 5'h18;
  assign when_Debug_l71_8 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_8_1);
  assign MulEU_MulEuPlugin_gprWritePort_valid = ((MulEU_MulEuPlugin_logicPhase_completesSuccessfully && MulEU_MulEuPlugin_euResult_writesToPreg) && (! MulEU_MulEuPlugin_euResult_destIsFpr));
  assign MulEU_MulEuPlugin_gprWritePort_address = MulEU_MulEuPlugin_euResult_uop_physDest_idx;
  assign MulEU_MulEuPlugin_gprWritePort_data = MulEU_MulEuPlugin_euResult_data;
  assign MulEU_MulEuPlugin_bypassOutputPort_valid = MulEU_MulEuPlugin_logicPhase_executionCompletes;
  assign MulEU_MulEuPlugin_bypassOutputPort_payload_physRegIdx = MulEU_MulEuPlugin_euResult_uop_physDest_idx;
  assign MulEU_MulEuPlugin_bypassOutputPort_payload_physRegData = MulEU_MulEuPlugin_euResult_data;
  assign MulEU_MulEuPlugin_bypassOutputPort_payload_robPtr = MulEU_MulEuPlugin_euResult_uop_robPtr;
  assign MulEU_MulEuPlugin_bypassOutputPort_payload_isFPR = MulEU_MulEuPlugin_euResult_destIsFpr;
  assign MulEU_MulEuPlugin_bypassOutputPort_payload_hasException = MulEU_MulEuPlugin_euResult_hasException;
  assign MulEU_MulEuPlugin_bypassOutputPort_payload_exceptionCode = MulEU_MulEuPlugin_euResult_exceptionCode;
  assign MulEU_MulEuPlugin_wakeupSourcePort_valid = (MulEU_MulEuPlugin_logicPhase_executionCompletes && MulEU_MulEuPlugin_euResult_writesToPreg);
  assign MulEU_MulEuPlugin_wakeupSourcePort_payload_physRegIdx = MulEU_MulEuPlugin_euResult_uop_physDest_idx;
  assign MulEU_MulEuPlugin_setup_clearBusyPort_valid = (MulEU_MulEuPlugin_logicPhase_executionCompletes && MulEU_MulEuPlugin_euResult_writesToPreg);
  assign MulEU_MulEuPlugin_setup_clearBusyPort_payload = MulEU_MulEuPlugin_euResult_uop_physDest_idx;
  assign when_EuBasePlugin_l300_1 = ((MulEU_MulEuPlugin_logicPhase_executionCompletes && MulEU_MulEuPlugin_euResult_writesToPreg) && (MulEU_MulEuPlugin_euResult_uop_physDest_idx < 6'h06));
  assign s0_Dispatch_valid_1 = BranchEU_BranchEuPlugin_euInputPort_valid;
  assign BranchEU_BranchEuPlugin_euInputPort_ready = s0_Dispatch_ready;
  assign _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3 = BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_condition;
  assign _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3 = BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_rtype;
  assign _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_3 = BranchEU_BranchEuPlugin_euInputPort_payload_pc;
  assign s0_Dispatch_isFiring = (s0_Dispatch_valid_1 && s0_Dispatch_ready);
  assign s1_Calc_isFiring = (s1_Calc_valid && s1_Calc_ready);
  assign BranchEU_BranchEuPlugin_gprReadPorts_0_valid = (s1_Calc_isFiring && _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_valid);
  assign BranchEU_BranchEuPlugin_gprReadPorts_0_address = _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_address;
  assign BranchEU_BranchEuPlugin_gprReadPorts_1_valid = (s1_Calc_isFiring && _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_valid);
  assign BranchEU_BranchEuPlugin_gprReadPorts_1_address = _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_address;
  always @(*) begin
    case(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2)
      BranchCondition_EQ : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = (BranchEU_BranchEuPlugin_gprReadPorts_0_rsp == BranchEU_BranchEuPlugin_gprReadPorts_1_rsp);
      end
      BranchCondition_NE : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = (BranchEU_BranchEuPlugin_gprReadPorts_0_rsp != BranchEU_BranchEuPlugin_gprReadPorts_1_rsp);
      end
      BranchCondition_LT : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = ($signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_3) < $signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_1));
      end
      BranchCondition_GE : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = ($signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_2) <= $signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_3));
      end
      BranchCondition_LTU : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = (BranchEU_BranchEuPlugin_gprReadPorts_0_rsp < BranchEU_BranchEuPlugin_gprReadPorts_1_rsp);
      end
      BranchCondition_GEU : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = (BranchEU_BranchEuPlugin_gprReadPorts_1_rsp <= BranchEU_BranchEuPlugin_gprReadPorts_0_rsp);
      end
      BranchCondition_EQZ : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = (BranchEU_BranchEuPlugin_gprReadPorts_0_rsp == 32'h0);
      end
      BranchCondition_NEZ : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = (BranchEU_BranchEuPlugin_gprReadPorts_0_rsp != 32'h0);
      end
      BranchCondition_LTZ : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = ($signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_4) < $signed(32'h0));
      end
      BranchCondition_GEZ : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = ($signed(32'h0) <= $signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_5));
      end
      BranchCondition_GTZ : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = ($signed(32'h0) < $signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_6));
      end
      BranchCondition_LEZ : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = ($signed(_zz__zz_BranchEU_BranchEuPlugin_euResult_data_3_7) <= $signed(32'h0));
      end
      default : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_3 = 1'b1;
      end
    endcase
  end

  assign switch_BranchEuPlugin_l133 = {_zz_switch_BranchEuPlugin_l133,_zz_switch_BranchEuPlugin_l133_1};
  always @(*) begin
    case(switch_BranchEuPlugin_l133)
      2'b00 : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_4 = (_zz_BranchEU_BranchEuPlugin_euResult_uop_pc_2 + _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4);
      end
      2'b01 : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_4 = _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_1;
      end
      2'b10 : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_4 = (_zz_BranchEU_BranchEuPlugin_euResult_uop_pc_2 + _zz__zz_BranchEU_BranchEuPlugin_euResult_data_4_4);
      end
      default : begin
        _zz_BranchEU_BranchEuPlugin_euResult_data_4 = (_zz_BranchEU_BranchEuPlugin_euResult_uop_pc_2 + 32'h00000004);
      end
    endcase
  end

  assign s2_Select_isFiring = (s2_Select_valid && s2_Select_ready);
  assign _zz_BranchEU_BranchEuPlugin_euResult_data_5 = (_zz_BranchEU_BranchEuPlugin_euResult_uop_pc_1 + 32'h00000004);
  always @(*) begin
    if(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump_1) begin
      _zz_BranchEU_BranchEuPlugin_euResult_isTaken_1 = 1'b1;
    end else begin
      _zz_BranchEU_BranchEuPlugin_euResult_isTaken_1 = _zz_BranchEU_BranchEuPlugin_euResult_data_2;
    end
  end

  always @(*) begin
    if(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump_1) begin
      _zz_BranchEU_BranchEuPlugin_euResult_data_6 = _zz_BranchEU_BranchEuPlugin_euResult_data_1;
    end else begin
      _zz_BranchEU_BranchEuPlugin_euResult_data_6 = (_zz_BranchEU_BranchEuPlugin_euResult_data_2 ? _zz_BranchEU_BranchEuPlugin_euResult_data_1 : _zz_BranchEU_BranchEuPlugin_euResult_data_5);
    end
  end

  always @(*) begin
    if(_zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted_1) begin
      _zz_BranchEU_BranchEuPlugin_euResult_isMispredictedBranch_1 = ((_zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken_1 == _zz_BranchEU_BranchEuPlugin_euResult_isTaken_1) && ((! _zz_BranchEU_BranchEuPlugin_euResult_isTaken_1) || (_zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target_1 == _zz_BranchEU_BranchEuPlugin_euResult_data_6)));
    end else begin
      _zz_BranchEU_BranchEuPlugin_euResult_isMispredictedBranch_1 = (! _zz_BranchEU_BranchEuPlugin_euResult_isTaken_1);
    end
  end

  assign _zz_52 = (! _zz_BranchEU_BranchEuPlugin_euResult_isMispredictedBranch_1);
  assign s3_Result_isFiring = (s3_Result_valid && s3_Result_ready);
  assign s3_Result_isFlushed = ROBPlugin_aggregatedFlushSignal_valid;
  assign when_Connection_l66_9 = (|{ROBPlugin_aggregatedFlushSignal_valid,ROBPlugin_aggregatedFlushSignal_valid});
  assign s2_Select_isFlushed = when_Connection_l66_9;
  assign when_Connection_l66_10 = (|{when_Connection_l66_9,ROBPlugin_aggregatedFlushSignal_valid});
  assign s1_Calc_isFlushed = when_Connection_l66_10;
  assign s0_Dispatch_isFlushed = (|{when_Connection_l66_10,ROBPlugin_aggregatedFlushSignal_valid});
  assign s0_Dispatch_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign s1_Calc_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign s2_Select_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  assign s3_Result_isFlushingRoot = (|ROBPlugin_aggregatedFlushSignal_valid);
  always @(*) begin
    _zz_s1_Calc_valid = s0_Dispatch_valid_1;
    if(s0_Dispatch_isFlushingRoot) begin
      _zz_s1_Calc_valid = 1'b0;
    end
  end

  assign s0_Dispatch_ready = 1'b1;
  always @(*) begin
    _zz_s2_Select_valid = s1_Calc_valid;
    if(s1_Calc_isFlushingRoot) begin
      _zz_s2_Select_valid = 1'b0;
    end
  end

  assign s1_Calc_ready = 1'b1;
  always @(*) begin
    _zz_s3_Result_valid = s2_Select_valid;
    if(s2_Select_isFlushingRoot) begin
      _zz_s3_Result_valid = 1'b0;
    end
  end

  assign s2_Select_ready = 1'b1;
  assign s3_Result_ready = 1'b1;
  assign when_EuBasePlugin_l230_2 = (ROBPlugin_aggregatedFlushSignal_valid && BranchEU_BranchEuPlugin_euResult_valid);
  assign BranchEU_BranchEuPlugin_logicPhase_executionCompletes = (BranchEU_BranchEuPlugin_euResult_valid && (! ROBPlugin_aggregatedFlushSignal_valid));
  assign BranchEU_BranchEuPlugin_logicPhase_completesSuccessfully = (BranchEU_BranchEuPlugin_logicPhase_executionCompletes && (! BranchEU_BranchEuPlugin_euResult_hasException));
  assign oneShot_23_io_triggerIn = (BranchEU_BranchEuPlugin_logicPhase_executionCompletes && (_zz_when_Debug_l71 < _zz_io_triggerIn_18));
  assign _zz_when_Debug_l71_10 = 5'h18;
  assign when_Debug_l71_9 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_9_1);
  assign BranchEU_BranchEuPlugin_gprWritePort_valid = ((BranchEU_BranchEuPlugin_logicPhase_completesSuccessfully && BranchEU_BranchEuPlugin_euResult_writesToPreg) && (! BranchEU_BranchEuPlugin_euResult_destIsFpr));
  assign BranchEU_BranchEuPlugin_gprWritePort_address = BranchEU_BranchEuPlugin_euResult_uop_physDest_idx;
  assign BranchEU_BranchEuPlugin_gprWritePort_data = BranchEU_BranchEuPlugin_euResult_data;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_valid = BranchEU_BranchEuPlugin_logicPhase_executionCompletes;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_payload_physRegIdx = BranchEU_BranchEuPlugin_euResult_uop_physDest_idx;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_payload_physRegData = BranchEU_BranchEuPlugin_euResult_data;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_payload_robPtr = BranchEU_BranchEuPlugin_euResult_uop_robPtr;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_payload_isFPR = BranchEU_BranchEuPlugin_euResult_destIsFpr;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_payload_hasException = BranchEU_BranchEuPlugin_euResult_hasException;
  assign BranchEU_BranchEuPlugin_bypassOutputPort_payload_exceptionCode = BranchEU_BranchEuPlugin_euResult_exceptionCode;
  assign BranchEU_BranchEuPlugin_wakeupSourcePort_valid = (BranchEU_BranchEuPlugin_logicPhase_executionCompletes && BranchEU_BranchEuPlugin_euResult_writesToPreg);
  assign BranchEU_BranchEuPlugin_wakeupSourcePort_payload_physRegIdx = BranchEU_BranchEuPlugin_euResult_uop_physDest_idx;
  assign BranchEU_BranchEuPlugin_setup_clearBusyPort_valid = (BranchEU_BranchEuPlugin_logicPhase_executionCompletes && BranchEU_BranchEuPlugin_euResult_writesToPreg);
  assign BranchEU_BranchEuPlugin_setup_clearBusyPort_payload = BranchEU_BranchEuPlugin_euResult_uop_physDest_idx;
  assign when_EuBasePlugin_l300_2 = ((BranchEU_BranchEuPlugin_logicPhase_executionCompletes && BranchEU_BranchEuPlugin_euResult_writesToPreg) && (BranchEU_BranchEuPlugin_euResult_uop_physDest_idx < 6'h06));
  assign LsuEU_LsuEuPlugin_hw_aguPort_flush = ROBPlugin_aggregatedFlushSignal_valid;
  assign _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize = LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_size;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_valid = LsuEU_LsuEuPlugin_euInputPort_valid;
  assign LsuEU_LsuEuPlugin_euInputPort_ready = LsuEU_LsuEuPlugin_euInputPort_translated_ready;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_qPtr = 3'b000;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_basePhysReg = LsuEU_LsuEuPlugin_euInputPort_payload_src1Tag;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_immediate = LsuEU_LsuEuPlugin_euInputPort_payload_imm;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize = _zz_LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_usePc = LsuEU_LsuEuPlugin_euInputPort_payload_usePc;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_pc = LsuEU_LsuEuPlugin_euInputPort_payload_pcData;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_dataReg = LsuEU_LsuEuPlugin_euInputPort_payload_src2Tag;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_robPtr = LsuEU_LsuEuPlugin_euInputPort_payload_robPtr;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_isLoad = (! LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isStore);
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_isStore = LsuEU_LsuEuPlugin_euInputPort_payload_memCtrl_isStore;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_isFlush = 1'b0;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_isIO = 1'b1;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_payload_physDst = LsuEU_LsuEuPlugin_euInputPort_payload_physDest_idx;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_valid = LsuEU_LsuEuPlugin_euInputPort_translated_valid;
  assign LsuEU_LsuEuPlugin_euInputPort_translated_ready = LsuEU_LsuEuPlugin_hw_aguPort_input_ready;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_qPtr = LsuEU_LsuEuPlugin_euInputPort_translated_payload_qPtr;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_basePhysReg = LsuEU_LsuEuPlugin_euInputPort_translated_payload_basePhysReg;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_immediate = LsuEU_LsuEuPlugin_euInputPort_translated_payload_immediate;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize = LsuEU_LsuEuPlugin_euInputPort_translated_payload_accessSize;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_usePc = LsuEU_LsuEuPlugin_euInputPort_translated_payload_usePc;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_pc = LsuEU_LsuEuPlugin_euInputPort_translated_payload_pc;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_dataReg = LsuEU_LsuEuPlugin_euInputPort_translated_payload_dataReg;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_robPtr = LsuEU_LsuEuPlugin_euInputPort_translated_payload_robPtr;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isLoad = LsuEU_LsuEuPlugin_euInputPort_translated_payload_isLoad;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isStore = LsuEU_LsuEuPlugin_euInputPort_translated_payload_isStore;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isFlush = LsuEU_LsuEuPlugin_euInputPort_translated_payload_isFlush;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isIO = LsuEU_LsuEuPlugin_euInputPort_translated_payload_isIO;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_payload_physDst = LsuEU_LsuEuPlugin_euInputPort_translated_payload_physDst;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_ready = streamDemux_1_io_input_ready;
  assign streamDemux_1_io_select = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isStore;
  assign io_outputs_0_combStage_valid = streamDemux_1_io_outputs_0_valid;
  assign io_outputs_0_combStage_payload_qPtr = streamDemux_1_io_outputs_0_payload_qPtr;
  assign io_outputs_0_combStage_payload_address = streamDemux_1_io_outputs_0_payload_address;
  assign io_outputs_0_combStage_payload_alignException = streamDemux_1_io_outputs_0_payload_alignException;
  assign io_outputs_0_combStage_payload_accessSize = streamDemux_1_io_outputs_0_payload_accessSize;
  assign io_outputs_0_combStage_payload_storeMask = streamDemux_1_io_outputs_0_payload_storeMask;
  assign io_outputs_0_combStage_payload_basePhysReg = streamDemux_1_io_outputs_0_payload_basePhysReg;
  assign io_outputs_0_combStage_payload_immediate = streamDemux_1_io_outputs_0_payload_immediate;
  assign io_outputs_0_combStage_payload_usePc = streamDemux_1_io_outputs_0_payload_usePc;
  assign io_outputs_0_combStage_payload_pc = streamDemux_1_io_outputs_0_payload_pc;
  assign io_outputs_0_combStage_payload_robPtr = streamDemux_1_io_outputs_0_payload_robPtr;
  assign io_outputs_0_combStage_payload_isLoad = streamDemux_1_io_outputs_0_payload_isLoad;
  assign io_outputs_0_combStage_payload_isStore = streamDemux_1_io_outputs_0_payload_isStore;
  assign io_outputs_0_combStage_payload_physDst = streamDemux_1_io_outputs_0_payload_physDst;
  assign io_outputs_0_combStage_payload_storeData = streamDemux_1_io_outputs_0_payload_storeData;
  assign io_outputs_0_combStage_payload_isFlush = streamDemux_1_io_outputs_0_payload_isFlush;
  assign io_outputs_0_combStage_payload_isIO = streamDemux_1_io_outputs_0_payload_isIO;
  assign io_outputs_1_combStage_valid = streamDemux_1_io_outputs_1_valid;
  assign io_outputs_1_combStage_payload_qPtr = streamDemux_1_io_outputs_1_payload_qPtr;
  assign io_outputs_1_combStage_payload_address = streamDemux_1_io_outputs_1_payload_address;
  assign io_outputs_1_combStage_payload_alignException = streamDemux_1_io_outputs_1_payload_alignException;
  assign io_outputs_1_combStage_payload_accessSize = streamDemux_1_io_outputs_1_payload_accessSize;
  assign io_outputs_1_combStage_payload_storeMask = streamDemux_1_io_outputs_1_payload_storeMask;
  assign io_outputs_1_combStage_payload_basePhysReg = streamDemux_1_io_outputs_1_payload_basePhysReg;
  assign io_outputs_1_combStage_payload_immediate = streamDemux_1_io_outputs_1_payload_immediate;
  assign io_outputs_1_combStage_payload_usePc = streamDemux_1_io_outputs_1_payload_usePc;
  assign io_outputs_1_combStage_payload_pc = streamDemux_1_io_outputs_1_payload_pc;
  assign io_outputs_1_combStage_payload_robPtr = streamDemux_1_io_outputs_1_payload_robPtr;
  assign io_outputs_1_combStage_payload_isLoad = streamDemux_1_io_outputs_1_payload_isLoad;
  assign io_outputs_1_combStage_payload_isStore = streamDemux_1_io_outputs_1_payload_isStore;
  assign io_outputs_1_combStage_payload_physDst = streamDemux_1_io_outputs_1_payload_physDst;
  assign io_outputs_1_combStage_payload_storeData = streamDemux_1_io_outputs_1_payload_storeData;
  assign io_outputs_1_combStage_payload_isFlush = streamDemux_1_io_outputs_1_payload_isFlush;
  assign io_outputs_1_combStage_payload_isIO = streamDemux_1_io_outputs_1_payload_isIO;
  assign _zz_io_outputs_0_combStage_translated_payload_size = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize;
  assign io_outputs_0_combStage_translated_valid = io_outputs_0_combStage_valid;
  assign io_outputs_0_combStage_ready = io_outputs_0_combStage_translated_ready;
  assign io_outputs_0_combStage_translated_payload_robPtr = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr;
  assign io_outputs_0_combStage_translated_payload_pdest = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst;
  assign io_outputs_0_combStage_translated_payload_address = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address;
  assign io_outputs_0_combStage_translated_payload_isIO = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO;
  assign io_outputs_0_combStage_translated_payload_size = _zz_io_outputs_0_combStage_translated_payload_size;
  assign io_outputs_0_combStage_translated_payload_hasEarlyException = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException;
  assign io_outputs_0_combStage_translated_payload_earlyExceptionCode = 8'h04;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_valid = io_outputs_0_combStage_translated_valid;
  assign io_outputs_0_combStage_translated_ready = LsuEU_LsuEuPlugin_hw_lqPushPort_ready;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_payload_robPtr = io_outputs_0_combStage_translated_payload_robPtr;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_payload_pdest = io_outputs_0_combStage_translated_payload_pdest;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_payload_address = io_outputs_0_combStage_translated_payload_address;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_payload_isIO = io_outputs_0_combStage_translated_payload_isIO;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_payload_size = io_outputs_0_combStage_translated_payload_size;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_payload_hasEarlyException = io_outputs_0_combStage_translated_payload_hasEarlyException;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_payload_earlyExceptionCode = io_outputs_0_combStage_translated_payload_earlyExceptionCode;
  assign _zz_io_outputs_1_combStage_translated_payload_accessSize = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize;
  assign io_outputs_1_combStage_translated_valid = io_outputs_1_combStage_valid;
  assign io_outputs_1_combStage_ready = io_outputs_1_combStage_translated_ready;
  assign io_outputs_1_combStage_translated_payload_addr = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address;
  assign io_outputs_1_combStage_translated_payload_data = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData;
  assign io_outputs_1_combStage_translated_payload_be = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask;
  assign io_outputs_1_combStage_translated_payload_robPtr = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr;
  assign io_outputs_1_combStage_translated_payload_accessSize = _zz_io_outputs_1_combStage_translated_payload_accessSize;
  assign io_outputs_1_combStage_translated_payload_isFlush = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush;
  assign io_outputs_1_combStage_translated_payload_isIO = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO;
  assign io_outputs_1_combStage_translated_payload_hasEarlyException = LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException;
  assign io_outputs_1_combStage_translated_payload_earlyExceptionCode = 8'h06;
  assign StoreBufferPlugin_hw_pushPortInst_valid = io_outputs_1_combStage_translated_valid;
  assign io_outputs_1_combStage_translated_ready = StoreBufferPlugin_hw_pushPortInst_ready;
  assign StoreBufferPlugin_hw_pushPortInst_payload_addr = io_outputs_1_combStage_translated_payload_addr;
  assign StoreBufferPlugin_hw_pushPortInst_payload_data = io_outputs_1_combStage_translated_payload_data;
  assign StoreBufferPlugin_hw_pushPortInst_payload_be = io_outputs_1_combStage_translated_payload_be;
  assign StoreBufferPlugin_hw_pushPortInst_payload_robPtr = io_outputs_1_combStage_translated_payload_robPtr;
  assign StoreBufferPlugin_hw_pushPortInst_payload_accessSize = io_outputs_1_combStage_translated_payload_accessSize;
  assign StoreBufferPlugin_hw_pushPortInst_payload_isFlush = io_outputs_1_combStage_translated_payload_isFlush;
  assign StoreBufferPlugin_hw_pushPortInst_payload_isIO = io_outputs_1_combStage_translated_payload_isIO;
  assign StoreBufferPlugin_hw_pushPortInst_payload_hasEarlyException = io_outputs_1_combStage_translated_payload_hasEarlyException;
  assign StoreBufferPlugin_hw_pushPortInst_payload_earlyExceptionCode = io_outputs_1_combStage_translated_payload_earlyExceptionCode;
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_fire = (LsuEU_LsuEuPlugin_hw_lqPushPort_valid && LsuEU_LsuEuPlugin_hw_lqPushPort_ready);
  assign StoreBufferPlugin_hw_pushPortInst_fire = (StoreBufferPlugin_hw_pushPortInst_valid && StoreBufferPlugin_hw_pushPortInst_ready);
  assign when_LsuEuPlugin_l141 = (LsuEU_LsuEuPlugin_hw_lqPushPort_fire || StoreBufferPlugin_hw_pushPortInst_fire);
  assign when_EuBasePlugin_l230_3 = (ROBPlugin_aggregatedFlushSignal_valid && LsuEU_LsuEuPlugin_euResult_valid);
  assign LsuEU_LsuEuPlugin_logicPhase_executionCompletes = (LsuEU_LsuEuPlugin_euResult_valid && (! ROBPlugin_aggregatedFlushSignal_valid));
  assign LsuEU_LsuEuPlugin_logicPhase_completesSuccessfully = (LsuEU_LsuEuPlugin_logicPhase_executionCompletes && (! LsuEU_LsuEuPlugin_euResult_hasException));
  assign oneShot_24_io_triggerIn = (LsuEU_LsuEuPlugin_logicPhase_executionCompletes && (_zz_when_Debug_l71 < _zz_io_triggerIn_20));
  assign _zz_when_Debug_l71_11 = 5'h18;
  assign when_Debug_l71_10 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_10_1);
  assign LsuEU_LsuEuPlugin_gprWritePort_valid = ((LsuEU_LsuEuPlugin_logicPhase_completesSuccessfully && LsuEU_LsuEuPlugin_euResult_writesToPreg) && (! LsuEU_LsuEuPlugin_euResult_destIsFpr));
  assign LsuEU_LsuEuPlugin_gprWritePort_address = LsuEU_LsuEuPlugin_euResult_uop_physDest_idx;
  assign LsuEU_LsuEuPlugin_gprWritePort_data = LsuEU_LsuEuPlugin_euResult_data;
  assign LsuEU_LsuEuPlugin_bypassOutputPort_valid = LsuEU_LsuEuPlugin_logicPhase_executionCompletes;
  assign LsuEU_LsuEuPlugin_bypassOutputPort_payload_physRegIdx = LsuEU_LsuEuPlugin_euResult_uop_physDest_idx;
  assign LsuEU_LsuEuPlugin_bypassOutputPort_payload_physRegData = LsuEU_LsuEuPlugin_euResult_data;
  assign LsuEU_LsuEuPlugin_bypassOutputPort_payload_robPtr = LsuEU_LsuEuPlugin_euResult_uop_robPtr;
  assign LsuEU_LsuEuPlugin_bypassOutputPort_payload_isFPR = LsuEU_LsuEuPlugin_euResult_destIsFpr;
  assign LsuEU_LsuEuPlugin_bypassOutputPort_payload_hasException = LsuEU_LsuEuPlugin_euResult_hasException;
  assign LsuEU_LsuEuPlugin_bypassOutputPort_payload_exceptionCode = LsuEU_LsuEuPlugin_euResult_exceptionCode;
  assign LsuEU_LsuEuPlugin_wakeupSourcePort_valid = (LsuEU_LsuEuPlugin_logicPhase_executionCompletes && LsuEU_LsuEuPlugin_euResult_writesToPreg);
  assign LsuEU_LsuEuPlugin_wakeupSourcePort_payload_physRegIdx = LsuEU_LsuEuPlugin_euResult_uop_physDest_idx;
  assign LsuEU_LsuEuPlugin_setup_clearBusyPort_valid = (LsuEU_LsuEuPlugin_logicPhase_executionCompletes && LsuEU_LsuEuPlugin_euResult_writesToPreg);
  assign LsuEU_LsuEuPlugin_setup_clearBusyPort_payload = LsuEU_LsuEuPlugin_euResult_uop_physDest_idx;
  assign when_EuBasePlugin_l300_3 = ((LsuEU_LsuEuPlugin_logicPhase_executionCompletes && LsuEU_LsuEuPlugin_euResult_writesToPreg) && (LsuEU_LsuEuPlugin_euResult_uop_physDest_idx < 6'h06));
  assign s3_Dispatch_isFlushed = when_Connection_l66;
  assign s2_RobAlloc_isFlushed = when_Connection_l66;
  assign when_Connection_l66_11 = (|{when_Connection_l66,_zz_s1_Rename_isFlushingRoot});
  assign s1_Rename_isFlushed = when_Connection_l66_11;
  assign s0_Decode_isFlushed = (|{when_Connection_l66_11,_zz_s0_Decode_isFlushingRoot});
  assign s0_Decode_isFlushingRoot = (|_zz_s0_Decode_isFlushingRoot);
  assign s1_Rename_isFlushingRoot = (|_zz_s1_Rename_isFlushingRoot);
  assign s3_Dispatch_isFlushingRoot = (|when_Connection_l66);
  always @(*) begin
    _zz_s1_Rename_valid = s0_Decode_valid;
    if(s0_Decode_isFlushingRoot) begin
      _zz_s1_Rename_valid = 1'b0;
    end
  end

  assign s0_Decode_ready = s0_Decode_ready_output;
  always @(*) begin
    _zz_s2_RobAlloc_valid = s1_Rename_valid;
    if(s1_Rename_isFlushingRoot) begin
      _zz_s2_RobAlloc_valid = 1'b0;
    end
  end

  assign s1_Rename_ready = s1_Rename_ready_output;
  always @(*) begin
    _zz_s3_Dispatch_valid = s2_RobAlloc_valid;
    if(when_Pipeline_l282) begin
      _zz_s3_Dispatch_valid = 1'b0;
    end
  end

  always @(*) begin
    s2_RobAlloc_ready = s2_RobAlloc_ready_output;
    if(when_Pipeline_l282) begin
      s2_RobAlloc_ready = 1'b0;
    end
  end

  assign when_Pipeline_l282 = (|{s2_RobAlloc_haltRequest_RobAllocPlugin_l30,s2_RobAlloc_haltRequest_RenamePlugin_l85});
  always @(*) begin
    s3_Dispatch_ready = 1'b1;
    if(when_Pipeline_l282_1) begin
      s3_Dispatch_ready = 1'b0;
    end
  end

  assign when_Pipeline_l282_1 = (|s3_Dispatch_haltRequest_DispatchPlugin_l78);
  always @(*) begin
    s0_Decode_ready_output = s1_Rename_ready;
    if(when_Connection_l74) begin
      s0_Decode_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74 = (! s1_Rename_valid);
  always @(*) begin
    s1_Rename_ready_output = s2_RobAlloc_ready;
    if(when_Connection_l74_1) begin
      s1_Rename_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_1 = (! s2_RobAlloc_valid);
  always @(*) begin
    s2_RobAlloc_ready_output = s3_Dispatch_ready;
    if(when_Connection_l74_2) begin
      s2_RobAlloc_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_2 = (! s3_Dispatch_valid);
  assign _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid = (LsuEU_LsuEuPlugin_hw_aguPort_input_valid && LsuEU_LsuEuPlugin_hw_aguPort_input_ready);
  assign LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid = _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid;
  assign LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_address = LsuEU_LsuEuPlugin_hw_aguPort_input_payload_basePhysReg;
  assign LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_valid = (_zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid && LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isStore);
  assign LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_address = LsuEU_LsuEuPlugin_hw_aguPort_input_payload_dataReg;
  always @(*) begin
    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_1 = 1'b0;
    if(AguPlugin_logic_bypassFlow_valid) begin
      if(when_AddressGenerationUnit_l215) begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_1 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_2 = 32'h0;
    if(AguPlugin_logic_bypassFlow_valid) begin
      if(when_AddressGenerationUnit_l215) begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_2 = AguPlugin_logic_bypassFlow_payload_physRegData;
      end
    end
  end

  always @(*) begin
    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_1 = 1'b0;
    if(AguPlugin_logic_bypassFlow_valid) begin
      if(when_AddressGenerationUnit_l220) begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_1 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_2 = 32'h0;
    if(AguPlugin_logic_bypassFlow_valid) begin
      if(when_AddressGenerationUnit_l220) begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_2 = AguPlugin_logic_bypassFlow_payload_physRegData;
      end
    end
  end

  assign when_AddressGenerationUnit_l215 = (AguPlugin_logic_bypassFlow_payload_physRegIdx == _zz_when_AddressGenerationUnit_l215);
  assign when_AddressGenerationUnit_l220 = (_zz_when_AddressGenerationUnit_l220_1 && (AguPlugin_logic_bypassFlow_payload_physRegIdx == _zz_when_AddressGenerationUnit_l220));
  assign _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_3 = (_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_1 ? _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_2 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address);
  always @(*) begin
    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_3 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(_zz_when_AddressGenerationUnit_l220_1) begin
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_3 = (_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_1 ? _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_2 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData);
    end
  end

  assign _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_4 = ((_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc ? _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc : _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_3) + _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate);
  always @(*) begin
    case(_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException)
      MemAccessSize_B : begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_1 = 3'b000;
      end
      MemAccessSize_H : begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_1 = 3'b001;
      end
      MemAccessSize_W : begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_1 = 3'b011;
      end
      default : begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_1 = 3'b111;
      end
    endcase
  end

  assign _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_4[1 : 0];
  always @(*) begin
    case(_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException)
      MemAccessSize_B : begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_1 = (4'b0001 <<< _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask);
      end
      MemAccessSize_H : begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_1 = (4'b0011 <<< (_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask & (~ 2'b01)));
      end
      MemAccessSize_W : begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_1 = 4'b1111;
      end
      default : begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_1 = 4'b1000;
      end
    endcase
  end

  assign _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException;
  always @(*) begin
    _zz_LsuEU_LsuEuPlugin_hw_aguPort_input_ready = LsuEU_LsuEuPlugin_hw_aguPort_output_ready;
    if(when_Stream_l477_5) begin
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_input_ready = 1'b1;
    end
  end

  assign when_Stream_l477_5 = (! _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid_1);
  assign _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid_1 = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid_2;
  assign _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1 = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_valid = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_5;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_2;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_2;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_basePhysReg = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_basePhysReg;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isStore = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isStore;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_4;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO = _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO_1;
  assign LsuEU_LsuEuPlugin_hw_aguPort_input_ready = (_zz_LsuEU_LsuEuPlugin_hw_aguPort_input_ready && (! LsuEU_LsuEuPlugin_hw_aguPort_flush));
  assign LsuEU_LsuEuPlugin_hw_lqPushPort_ready = streamArbiter_9_io_inputs_0_ready;
  assign LoadQueuePlugin_logic_pushCmd_valid = streamArbiter_9_io_output_valid;
  assign LoadQueuePlugin_logic_pushCmd_payload_robPtr = streamArbiter_9_io_output_payload_robPtr;
  assign LoadQueuePlugin_logic_pushCmd_payload_pdest = streamArbiter_9_io_output_payload_pdest;
  assign LoadQueuePlugin_logic_pushCmd_payload_address = streamArbiter_9_io_output_payload_address;
  assign LoadQueuePlugin_logic_pushCmd_payload_isIO = streamArbiter_9_io_output_payload_isIO;
  assign LoadQueuePlugin_logic_pushCmd_payload_size = streamArbiter_9_io_output_payload_size;
  assign LoadQueuePlugin_logic_pushCmd_payload_hasEarlyException = streamArbiter_9_io_output_payload_hasEarlyException;
  assign LoadQueuePlugin_logic_pushCmd_payload_earlyExceptionCode = streamArbiter_9_io_output_payload_earlyExceptionCode;
  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_completionInfo_valid = 1'b0;
    if(LoadQueuePlugin_logic_loadQueue_popOnFwdHit) begin
      LoadQueuePlugin_logic_loadQueue_completionInfo_valid = 1'b1;
    end else begin
      if(LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess) begin
        LoadQueuePlugin_logic_loadQueue_completionInfo_valid = 1'b1;
      end else begin
        if(LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead) begin
          LoadQueuePlugin_logic_loadQueue_completionInfo_valid = 1'b1;
        end else begin
          if(LoadQueuePlugin_logic_loadQueue_popOnEarlyException) begin
            LoadQueuePlugin_logic_loadQueue_completionInfo_valid = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_completionInfo_fromFwd = 1'b0;
    if(LoadQueuePlugin_logic_loadQueue_popOnFwdHit) begin
      LoadQueuePlugin_logic_loadQueue_completionInfo_fromFwd = 1'b1;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_completionInfo_fromDCache = 1'b0;
    if(!LoadQueuePlugin_logic_loadQueue_popOnFwdHit) begin
      if(LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess) begin
        LoadQueuePlugin_logic_loadQueue_completionInfo_fromDCache = 1'b1;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_completionInfo_fromMMIO = 1'b0;
    if(!LoadQueuePlugin_logic_loadQueue_popOnFwdHit) begin
      if(!LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess) begin
        if(LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead) begin
          LoadQueuePlugin_logic_loadQueue_completionInfo_fromMMIO = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_completionInfo_fromEarlyExc = 1'b0;
    if(!LoadQueuePlugin_logic_loadQueue_popOnFwdHit) begin
      if(!LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess) begin
        if(!LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead) begin
          if(LoadQueuePlugin_logic_loadQueue_popOnEarlyException) begin
            LoadQueuePlugin_logic_loadQueue_completionInfo_fromEarlyExc = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_completionInfo_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(LoadQueuePlugin_logic_loadQueue_popOnFwdHit) begin
      LoadQueuePlugin_logic_loadQueue_completionInfo_data = LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_data;
    end else begin
      if(LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess) begin
        LoadQueuePlugin_logic_loadQueue_completionInfo_data = LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_data;
      end else begin
        if(LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead) begin
          LoadQueuePlugin_logic_loadQueue_completionInfo_data = CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_payload_data;
        end
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_completionInfo_hasFault = 1'b0;
    if(LoadQueuePlugin_logic_loadQueue_popOnFwdHit) begin
      LoadQueuePlugin_logic_loadQueue_completionInfo_hasFault = 1'b0;
    end else begin
      if(LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess) begin
        LoadQueuePlugin_logic_loadQueue_completionInfo_hasFault = LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_fault;
      end else begin
        if(LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead) begin
          LoadQueuePlugin_logic_loadQueue_completionInfo_hasFault = CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_payload_error;
        end else begin
          if(LoadQueuePlugin_logic_loadQueue_popOnEarlyException) begin
            LoadQueuePlugin_logic_loadQueue_completionInfo_hasFault = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_completionInfo_exceptionCode = 8'bxxxxxxxx;
    if(!LoadQueuePlugin_logic_loadQueue_popOnFwdHit) begin
      if(LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess) begin
        LoadQueuePlugin_logic_loadQueue_completionInfo_exceptionCode = 8'h05;
      end else begin
        if(LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead) begin
          LoadQueuePlugin_logic_loadQueue_completionInfo_exceptionCode = 8'h05;
        end else begin
          if(LoadQueuePlugin_logic_loadQueue_popOnEarlyException) begin
            LoadQueuePlugin_logic_loadQueue_completionInfo_exceptionCode = LoadQueuePlugin_logic_loadQueue_slots_0_exceptionCode;
          end
        end
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_valid = LoadQueuePlugin_logic_loadQueue_slots_0_valid;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_address = LoadQueuePlugin_logic_loadQueue_slots_0_address;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_address = LoadQueuePlugin_logic_pushCmd_payload_address;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size = LoadQueuePlugin_logic_loadQueue_slots_0_size;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size = LoadQueuePlugin_logic_pushCmd_payload_size;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_robPtr = LoadQueuePlugin_logic_loadQueue_slots_0_robPtr;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_robPtr = LoadQueuePlugin_logic_pushCmd_payload_robPtr;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_pdest = LoadQueuePlugin_logic_loadQueue_slots_0_pdest;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_pdest = LoadQueuePlugin_logic_pushCmd_payload_pdest;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isIO = LoadQueuePlugin_logic_loadQueue_slots_0_isIO;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isIO = LoadQueuePlugin_logic_pushCmd_payload_isIO;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_hasException = LoadQueuePlugin_logic_loadQueue_slots_0_hasException;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_hasException = LoadQueuePlugin_logic_pushCmd_payload_hasEarlyException;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_exceptionCode = LoadQueuePlugin_logic_loadQueue_slots_0_exceptionCode;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_exceptionCode = LoadQueuePlugin_logic_pushCmd_payload_earlyExceptionCode;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForFwdRsp = 1'b0;
      end
    end
    if(StoreBufferPlugin_hw_sqQueryPort_cmd_valid) begin
      LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForFwdRsp = 1'b1;
    end
    if(when_LoadQueuePlugin_l329) begin
      LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForFwdRsp = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slots_0_isStalledByDependency;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isStalledByDependency = 1'b0;
      end
    end
    if(when_LoadQueuePlugin_l329) begin
      if(!LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_hit) begin
        if(when_LoadQueuePlugin_l335) begin
          LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isStalledByDependency = 1'b1;
        end
      end
    end
    if(LoadQueuePlugin_logic_loadQueue_slots_0_isStalledByDependency) begin
      LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isStalledByDependency = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache = 1'b0;
      end
    end
    if(when_LoadQueuePlugin_l329) begin
      if(!LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_hit) begin
        if(!when_LoadQueuePlugin_l335) begin
          LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache = 1'b1;
        end
      end
    end
    if(when_LoadQueuePlugin_l350) begin
      LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache = 1'b1;
    end
    if(LoadQueuePlugin_hw_dCacheLoadPort_cmd_fire) begin
      LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_mmioCmdFired) begin
      LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache = 1'b0;
    end
    if(when_LoadQueuePlugin_l409) begin
      if(LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_redo) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache = 1'b1;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_54) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForRsp = 1'b0;
      end
    end
    if(LoadQueuePlugin_hw_dCacheLoadPort_cmd_fire) begin
      LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForRsp = 1'b1;
    end
    if(LoadQueuePlugin_logic_loadQueue_mmioCmdFired) begin
      LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForRsp = 1'b1;
    end
    if(when_LoadQueuePlugin_l409) begin
      if(LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_redo) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForRsp = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_valid = LoadQueuePlugin_logic_loadQueue_slots_1_valid;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_address = LoadQueuePlugin_logic_loadQueue_slots_1_address;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_address = LoadQueuePlugin_logic_pushCmd_payload_address;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size = LoadQueuePlugin_logic_loadQueue_slots_1_size;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size = LoadQueuePlugin_logic_pushCmd_payload_size;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_robPtr = LoadQueuePlugin_logic_loadQueue_slots_1_robPtr;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_robPtr = LoadQueuePlugin_logic_pushCmd_payload_robPtr;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_pdest = LoadQueuePlugin_logic_loadQueue_slots_1_pdest;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_pdest = LoadQueuePlugin_logic_pushCmd_payload_pdest;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isIO = LoadQueuePlugin_logic_loadQueue_slots_1_isIO;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isIO = LoadQueuePlugin_logic_pushCmd_payload_isIO;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_hasException = LoadQueuePlugin_logic_loadQueue_slots_1_hasException;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_hasException = LoadQueuePlugin_logic_pushCmd_payload_hasEarlyException;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_exceptionCode = LoadQueuePlugin_logic_loadQueue_slots_1_exceptionCode;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_exceptionCode = LoadQueuePlugin_logic_pushCmd_payload_earlyExceptionCode;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slots_1_isWaitingForFwdRsp;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForFwdRsp = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slots_1_isStalledByDependency;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isStalledByDependency = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slots_1_isReadyForDCache;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isReadyForDCache = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slots_1_isWaitingForRsp;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_55) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForRsp = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_valid = LoadQueuePlugin_logic_loadQueue_slots_2_valid;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_address = LoadQueuePlugin_logic_loadQueue_slots_2_address;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_address = LoadQueuePlugin_logic_pushCmd_payload_address;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size = LoadQueuePlugin_logic_loadQueue_slots_2_size;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size = LoadQueuePlugin_logic_pushCmd_payload_size;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_robPtr = LoadQueuePlugin_logic_loadQueue_slots_2_robPtr;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_robPtr = LoadQueuePlugin_logic_pushCmd_payload_robPtr;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_pdest = LoadQueuePlugin_logic_loadQueue_slots_2_pdest;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_pdest = LoadQueuePlugin_logic_pushCmd_payload_pdest;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isIO = LoadQueuePlugin_logic_loadQueue_slots_2_isIO;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isIO = LoadQueuePlugin_logic_pushCmd_payload_isIO;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_hasException = LoadQueuePlugin_logic_loadQueue_slots_2_hasException;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_hasException = LoadQueuePlugin_logic_pushCmd_payload_hasEarlyException;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_exceptionCode = LoadQueuePlugin_logic_loadQueue_slots_2_exceptionCode;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_exceptionCode = LoadQueuePlugin_logic_pushCmd_payload_earlyExceptionCode;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slots_2_isWaitingForFwdRsp;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForFwdRsp = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slots_2_isStalledByDependency;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isStalledByDependency = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slots_2_isReadyForDCache;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isReadyForDCache = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slots_2_isWaitingForRsp;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_56) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForRsp = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_valid = LoadQueuePlugin_logic_loadQueue_slots_3_valid;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_address = LoadQueuePlugin_logic_loadQueue_slots_3_address;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_address = LoadQueuePlugin_logic_pushCmd_payload_address;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size = LoadQueuePlugin_logic_loadQueue_slots_3_size;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size = LoadQueuePlugin_logic_pushCmd_payload_size;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_robPtr = LoadQueuePlugin_logic_loadQueue_slots_3_robPtr;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_robPtr = LoadQueuePlugin_logic_pushCmd_payload_robPtr;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_pdest = LoadQueuePlugin_logic_loadQueue_slots_3_pdest;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_pdest = LoadQueuePlugin_logic_pushCmd_payload_pdest;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isIO = LoadQueuePlugin_logic_loadQueue_slots_3_isIO;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isIO = LoadQueuePlugin_logic_pushCmd_payload_isIO;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_hasException = LoadQueuePlugin_logic_loadQueue_slots_3_hasException;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_hasException = LoadQueuePlugin_logic_pushCmd_payload_hasEarlyException;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_exceptionCode = LoadQueuePlugin_logic_loadQueue_slots_3_exceptionCode;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_exceptionCode = LoadQueuePlugin_logic_pushCmd_payload_earlyExceptionCode;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slots_3_isWaitingForFwdRsp;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForFwdRsp = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slots_3_isStalledByDependency;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isStalledByDependency = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slots_3_isReadyForDCache;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isReadyForDCache = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slots_3_isWaitingForRsp;
    if(LoadQueuePlugin_logic_pushCmd_fire) begin
      if(_zz_57) begin
        LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForRsp = 1'b0;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_valid = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_valid;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_valid = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_valid = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_valid;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_valid = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_address = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_address;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_address = 32'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_address = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_address;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_address = 32'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_size = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_size;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_size = MemAccessSize_W;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_size = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_size = MemAccessSize_W;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_robPtr = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_robPtr;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_robPtr = 4'b0000;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_robPtr = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_robPtr;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_pdest = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_pdest;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_pdest = 6'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_pdest = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_pdest;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_pdest = 6'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_isIO = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isIO;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isIO = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isIO = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isIO;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isIO = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_hasException = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_hasException;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_hasException = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_hasException = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_hasException;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_hasException = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_exceptionCode = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_exceptionCode;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_exceptionCode = 8'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_exceptionCode = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_exceptionCode;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_exceptionCode = 8'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForFwdRsp;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForFwdRsp = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForFwdRsp;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForFwdRsp = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isStalledByDependency;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isStalledByDependency = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isStalledByDependency;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isStalledByDependency = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isReadyForDCache;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isReadyForDCache = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isReadyForDCache;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isReadyForDCache = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_0_isWaitingForRsp;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForRsp = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForRsp;
    end
    if(when_LoadQueuePlugin_l508) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForRsp = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_valid = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_valid;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_valid = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_valid = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_valid;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_valid = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_address = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_address;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_address = 32'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_address = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_address;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_address = 32'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_size = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_size;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_size = MemAccessSize_W;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_size = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_size = MemAccessSize_W;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_robPtr = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_robPtr;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_robPtr = 4'b0000;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_robPtr = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_robPtr;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_pdest = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_pdest;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_pdest = 6'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_pdest = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_pdest;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_pdest = 6'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_isIO = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isIO;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isIO = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isIO = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isIO;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isIO = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_hasException = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_hasException;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_hasException = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_hasException = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_hasException;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_hasException = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_exceptionCode = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_exceptionCode;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_exceptionCode = 8'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_exceptionCode = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_exceptionCode;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_exceptionCode = 8'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForFwdRsp;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForFwdRsp = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForFwdRsp;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForFwdRsp = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isStalledByDependency;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isStalledByDependency = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isStalledByDependency;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isStalledByDependency = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isReadyForDCache;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isReadyForDCache = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isReadyForDCache;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isReadyForDCache = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_1_isWaitingForRsp;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForRsp = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForRsp;
    end
    if(when_LoadQueuePlugin_l508_1) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForRsp = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_valid = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_valid;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_valid = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_valid = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_valid;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_valid = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_address = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_address;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_address = 32'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_address = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_address;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_address = 32'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_size = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_size;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_size = MemAccessSize_W;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_size = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_size = MemAccessSize_W;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_robPtr = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_robPtr;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_robPtr = 4'b0000;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_robPtr = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_robPtr;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_pdest = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_pdest;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_pdest = 6'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_pdest = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_pdest;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_pdest = 6'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_isIO = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isIO;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isIO = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isIO = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isIO;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isIO = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_hasException = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_hasException;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_hasException = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_hasException = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_hasException;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_hasException = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_exceptionCode = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_exceptionCode;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_exceptionCode = 8'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_exceptionCode = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_exceptionCode;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_exceptionCode = 8'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForFwdRsp;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForFwdRsp = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForFwdRsp;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForFwdRsp = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isStalledByDependency;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isStalledByDependency = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isStalledByDependency;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isStalledByDependency = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isReadyForDCache;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isReadyForDCache = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isReadyForDCache;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isReadyForDCache = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_2_isWaitingForRsp;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForRsp = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForRsp;
    end
    if(when_LoadQueuePlugin_l508_2) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForRsp = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_valid = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_valid;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_valid = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_valid = 1'b0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_valid = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_address = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_address;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_address = 32'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_address = 32'h0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_address = 32'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_size = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_size;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_size = MemAccessSize_W;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_size = MemAccessSize_W;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_size = MemAccessSize_W;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_robPtr = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_robPtr;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_robPtr = 4'b0000;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_robPtr = 4'b0000;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_pdest = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_pdest;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_pdest = 6'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_pdest = 6'h0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_pdest = 6'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_isIO = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isIO;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isIO = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isIO = 1'b0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isIO = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_hasException = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_hasException;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_hasException = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_hasException = 1'b0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_hasException = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_exceptionCode = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_exceptionCode;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_exceptionCode = 8'h0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_exceptionCode = 8'h0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_exceptionCode = 8'h0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForFwdRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForFwdRsp;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForFwdRsp = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForFwdRsp = 1'b0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForFwdRsp = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_isStalledByDependency = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isStalledByDependency;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isStalledByDependency = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isStalledByDependency = 1'b0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isStalledByDependency = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_isReadyForDCache = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isReadyForDCache;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isReadyForDCache = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isReadyForDCache = 1'b0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isReadyForDCache = 1'b0;
    end
  end

  always @(*) begin
    LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForRsp = LoadQueuePlugin_logic_loadQueue_slotsAfterUpdates_3_isWaitingForRsp;
    if(when_LoadQueuePlugin_l291) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForRsp = 1'b0;
    end
    if(LoadQueuePlugin_logic_loadQueue_popRequest) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForRsp = 1'b0;
    end
    if(when_LoadQueuePlugin_l508_3) begin
      LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForRsp = 1'b0;
    end
  end

  assign LoadQueuePlugin_logic_loadQueue_flushInProgress = (ROBPlugin_aggregatedFlushSignal_valid && (ROBPlugin_aggregatedFlushSignal_payload_reason == FlushReason_ROLLBACK_TO_ROB_IDX));
  assign when_LoadQueuePlugin_l291 = (ROBPlugin_aggregatedFlushSignal_valid && (ROBPlugin_aggregatedFlushSignal_payload_reason == FlushReason_FULL_FLUSH));
  assign LoadQueuePlugin_logic_loadQueue_canPush = ((! (&{LoadQueuePlugin_logic_loadQueue_slots_3_valid,{LoadQueuePlugin_logic_loadQueue_slots_2_valid,{LoadQueuePlugin_logic_loadQueue_slots_1_valid,LoadQueuePlugin_logic_loadQueue_slots_0_valid}}})) && (! LoadQueuePlugin_logic_loadQueue_flushInProgress));
  assign LoadQueuePlugin_logic_pushCmd_ready = LoadQueuePlugin_logic_loadQueue_canPush;
  assign LoadQueuePlugin_logic_loadQueue_availableSlotsMask = {(! LoadQueuePlugin_logic_loadQueue_slots_3_valid),{(! LoadQueuePlugin_logic_loadQueue_slots_2_valid),{(! LoadQueuePlugin_logic_loadQueue_slots_1_valid),(! LoadQueuePlugin_logic_loadQueue_slots_0_valid)}}};
  assign LoadQueuePlugin_logic_loadQueue_pushOh = (LoadQueuePlugin_logic_loadQueue_availableSlotsMask & _zz_LoadQueuePlugin_logic_loadQueue_pushOh);
  assign _zz_LoadQueuePlugin_logic_loadQueue_pushIdx = LoadQueuePlugin_logic_loadQueue_pushOh[3];
  assign _zz_LoadQueuePlugin_logic_loadQueue_pushIdx_1 = (LoadQueuePlugin_logic_loadQueue_pushOh[1] || _zz_LoadQueuePlugin_logic_loadQueue_pushIdx);
  assign _zz_LoadQueuePlugin_logic_loadQueue_pushIdx_2 = (LoadQueuePlugin_logic_loadQueue_pushOh[2] || _zz_LoadQueuePlugin_logic_loadQueue_pushIdx);
  assign LoadQueuePlugin_logic_loadQueue_pushIdx = {_zz_LoadQueuePlugin_logic_loadQueue_pushIdx_2,_zz_LoadQueuePlugin_logic_loadQueue_pushIdx_1};
  assign LoadQueuePlugin_logic_pushCmd_fire = (LoadQueuePlugin_logic_pushCmd_valid && LoadQueuePlugin_logic_pushCmd_ready);
  assign _zz_53 = ({3'd0,1'b1} <<< LoadQueuePlugin_logic_loadQueue_pushIdx);
  assign _zz_54 = _zz_53[0];
  assign _zz_55 = _zz_53[1];
  assign _zz_56 = _zz_53[2];
  assign _zz_57 = _zz_53[3];
  assign _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible = LoadQueuePlugin_logic_loadQueue_slots_0_robPtr[3];
  assign _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_1 = LoadQueuePlugin_logic_loadQueue_slots_0_robPtr[2 : 0];
  assign _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_2 = ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr[3];
  assign _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_3 = ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr[2 : 0];
  assign LoadQueuePlugin_logic_loadQueue_headIsVisible = (LoadQueuePlugin_logic_loadQueue_slots_0_valid && (! (LoadQueuePlugin_logic_loadQueue_flushInProgress && (((_zz_LoadQueuePlugin_logic_loadQueue_headIsVisible == _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_2) && (_zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_3 <= _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_1)) || ((_zz_LoadQueuePlugin_logic_loadQueue_headIsVisible != _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_2) && (_zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_1 < _zz_LoadQueuePlugin_logic_loadQueue_headIsVisible_3))))));
  assign LoadQueuePlugin_logic_loadQueue_headIsReadyForFwdQuery = (((((LoadQueuePlugin_logic_loadQueue_headIsVisible && (! LoadQueuePlugin_logic_loadQueue_slots_0_hasException)) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp)) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isStalledByDependency)) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp)) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache));
  assign StoreBufferPlugin_hw_sqQueryPort_cmd_valid = LoadQueuePlugin_logic_loadQueue_headIsReadyForFwdQuery;
  assign StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address = LoadQueuePlugin_logic_loadQueue_slots_0_address;
  assign StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size = LoadQueuePlugin_logic_loadQueue_slots_0_size;
  assign StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr = LoadQueuePlugin_logic_loadQueue_slots_0_robPtr;
  assign when_LoadQueuePlugin_l329 = (LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp && LoadQueuePlugin_logic_loadQueue_sbQueryRspValid);
  assign when_LoadQueuePlugin_l335 = (LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_olderStoreHasUnknownAddress || LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_olderStoreDataNotReady);
  assign when_LoadQueuePlugin_l350 = ((((LoadQueuePlugin_logic_loadQueue_headIsVisible && LoadQueuePlugin_logic_loadQueue_slots_0_hasException) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache)) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp)) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp));
  assign LoadQueuePlugin_logic_loadQueue_headIsReadyToExecute = ((LoadQueuePlugin_logic_loadQueue_headIsVisible && LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp));
  assign LoadQueuePlugin_logic_loadQueue_shouldNotSendToMemory = (LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp || (LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp && StoreBufferPlugin_hw_sqQueryPort_rsp_hit));
  assign LoadQueuePlugin_hw_dCacheLoadPort_cmd_valid = (((LoadQueuePlugin_logic_loadQueue_headIsReadyToExecute && (! LoadQueuePlugin_logic_loadQueue_slots_0_hasException)) && (! LoadQueuePlugin_logic_loadQueue_shouldNotSendToMemory)) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isIO));
  assign LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_virtual = LoadQueuePlugin_logic_loadQueue_slots_0_address;
  always @(*) begin
    _zz_LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size = 2'b00;
    case(LoadQueuePlugin_logic_loadQueue_slots_0_size)
      MemAccessSize_B : begin
        _zz_LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size = 2'b00;
      end
      MemAccessSize_H : begin
        _zz_LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size = 2'b01;
      end
      MemAccessSize_W : begin
        _zz_LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size = 2'b10;
      end
      default : begin
        _zz_LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size = 2'b11;
      end
    endcase
  end

  assign LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size = _zz_LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_size;
  assign LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_redoOnDataHazard = 1'b1;
  assign LoadQueuePlugin_hw_dCacheLoadPort_cmd_payload_id = LoadQueuePlugin_logic_loadQueue_slots_0_robPtr[2:0];
  assign LoadQueuePlugin_hw_dCacheLoadPort_translated_physical = LoadQueuePlugin_logic_loadQueue_slots_0_address;
  assign LoadQueuePlugin_hw_dCacheLoadPort_translated_abord = LoadQueuePlugin_logic_loadQueue_slots_0_hasException;
  assign LoadQueuePlugin_hw_dCacheLoadPort_cancels = 3'b000;
  assign LoadQueuePlugin_hw_dCacheLoadPort_cmd_fire = (LoadQueuePlugin_hw_dCacheLoadPort_cmd_valid && LoadQueuePlugin_hw_dCacheLoadPort_cmd_ready);
  assign _zz_LoadQueuePlugin_logic_loadQueue_mmioCmdFired = (((LoadQueuePlugin_logic_loadQueue_headIsReadyToExecute && (! LoadQueuePlugin_logic_loadQueue_slots_0_hasException)) && (! LoadQueuePlugin_logic_loadQueue_shouldNotSendToMemory)) && LoadQueuePlugin_logic_loadQueue_slots_0_isIO);
  assign LoadQueuePlugin_logic_loadQueue_mmioCmdFired = (_zz_LoadQueuePlugin_logic_loadQueue_mmioCmdFired && CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_cmd_ready);
  assign LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead = (((CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_valid && LoadQueuePlugin_logic_loadQueue_slots_0_valid) && (LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp || LoadQueuePlugin_logic_loadQueue_mmioCmdFired)) && LoadQueuePlugin_logic_loadQueue_slots_0_isIO);
  assign when_LoadQueuePlugin_l409 = (((LoadQueuePlugin_hw_dCacheLoadPort_rsp_valid && LoadQueuePlugin_logic_loadQueue_slots_0_valid) && LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isIO));
  assign LoadQueuePlugin_logic_loadQueue_popOnFwdHit = (LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp && LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_hit);
  assign LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess = ((((LoadQueuePlugin_hw_dCacheLoadPort_rsp_valid && LoadQueuePlugin_logic_loadQueue_slots_0_valid) && LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isIO)) && (! LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_redo));
  assign LoadQueuePlugin_logic_loadQueue_popOnEarlyException = ((LoadQueuePlugin_logic_loadQueue_slots_0_valid && LoadQueuePlugin_logic_loadQueue_slots_0_hasException) && (! LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache));
  assign LoadQueuePlugin_logic_loadQueue_popRequest = (((LoadQueuePlugin_logic_loadQueue_popOnFwdHit || LoadQueuePlugin_logic_loadQueue_popOnDCacheSuccess) || LoadQueuePlugin_logic_loadQueue_mmioResponseIsForHead) || LoadQueuePlugin_logic_loadQueue_popOnEarlyException);
  always @(*) begin
    ROBPlugin_robComponent_io_writeback_4_fire = 1'b0;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      ROBPlugin_robComponent_io_writeback_4_fire = 1'b1;
    end
  end

  always @(*) begin
    ROBPlugin_robComponent_io_writeback_4_robPtr = 4'bxxxx;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      ROBPlugin_robComponent_io_writeback_4_robPtr = LoadQueuePlugin_logic_loadQueue_completingHead_robPtr;
    end
  end

  always @(*) begin
    ROBPlugin_robComponent_io_writeback_4_result = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      ROBPlugin_robComponent_io_writeback_4_result = LoadQueuePlugin_logic_loadQueue_completionInfoReg_data;
    end
  end

  always @(*) begin
    ROBPlugin_robComponent_io_writeback_4_exceptionOccurred = 1'bx;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      ROBPlugin_robComponent_io_writeback_4_exceptionOccurred = LoadQueuePlugin_logic_loadQueue_completionInfoReg_hasFault;
    end
  end

  always @(*) begin
    ROBPlugin_robComponent_io_writeback_4_exceptionCodeIn = 8'bxxxxxxxx;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      ROBPlugin_robComponent_io_writeback_4_exceptionCodeIn = LoadQueuePlugin_logic_loadQueue_completionInfoReg_exceptionCode;
    end
  end

  always @(*) begin
    LoadQueuePlugin_hw_prfWritePort_valid = 1'b0;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      if(when_LoadQueuePlugin_l478) begin
        LoadQueuePlugin_hw_prfWritePort_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_hw_prfWritePort_address = 6'bxxxxxx;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      if(when_LoadQueuePlugin_l478) begin
        LoadQueuePlugin_hw_prfWritePort_address = LoadQueuePlugin_logic_loadQueue_completingHead_pdest;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_hw_prfWritePort_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      if(when_LoadQueuePlugin_l478) begin
        LoadQueuePlugin_hw_prfWritePort_data = LoadQueuePlugin_logic_loadQueue_completionInfoReg_data;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_hw_wakeupPort_valid = 1'b0;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      if(when_LoadQueuePlugin_l478) begin
        LoadQueuePlugin_hw_wakeupPort_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_hw_wakeupPort_payload_physRegIdx = 6'bxxxxxx;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      if(when_LoadQueuePlugin_l478) begin
        LoadQueuePlugin_hw_wakeupPort_payload_physRegIdx = LoadQueuePlugin_logic_loadQueue_completingHead_pdest;
      end
    end
  end

  always @(*) begin
    LoadQueuePlugin_hw_busyTableClearPort_valid = 1'b0;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      LoadQueuePlugin_hw_busyTableClearPort_valid = 1'b1;
    end
  end

  always @(*) begin
    LoadQueuePlugin_hw_busyTableClearPort_payload = 6'bxxxxxx;
    if(LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid) begin
      LoadQueuePlugin_hw_busyTableClearPort_payload = LoadQueuePlugin_logic_loadQueue_completingHead_pdest;
    end
  end

  assign when_LoadQueuePlugin_l478 = (! LoadQueuePlugin_logic_loadQueue_completionInfoReg_hasFault);
  assign _zz_when_LoadQueuePlugin_l508 = LoadQueuePlugin_logic_loadQueue_slots_0_robPtr[3];
  assign _zz_when_LoadQueuePlugin_l508_1 = LoadQueuePlugin_logic_loadQueue_slots_0_robPtr[2 : 0];
  assign _zz_when_LoadQueuePlugin_l508_2 = LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr[3];
  assign _zz_when_LoadQueuePlugin_l508_3 = LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr[2 : 0];
  assign when_LoadQueuePlugin_l508 = ((LoadQueuePlugin_logic_loadQueue_registeredFlush_valid && LoadQueuePlugin_logic_loadQueue_slots_0_valid) && (((_zz_when_LoadQueuePlugin_l508 == _zz_when_LoadQueuePlugin_l508_2) && (_zz_when_LoadQueuePlugin_l508_3 <= _zz_when_LoadQueuePlugin_l508_1)) || ((_zz_when_LoadQueuePlugin_l508 != _zz_when_LoadQueuePlugin_l508_2) && (_zz_when_LoadQueuePlugin_l508_1 < _zz_when_LoadQueuePlugin_l508_3))));
  assign _zz_when_LoadQueuePlugin_l508_4 = LoadQueuePlugin_logic_loadQueue_slots_1_robPtr[3];
  assign _zz_when_LoadQueuePlugin_l508_5 = LoadQueuePlugin_logic_loadQueue_slots_1_robPtr[2 : 0];
  assign _zz_when_LoadQueuePlugin_l508_6 = LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr[3];
  assign _zz_when_LoadQueuePlugin_l508_7 = LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr[2 : 0];
  assign when_LoadQueuePlugin_l508_1 = ((LoadQueuePlugin_logic_loadQueue_registeredFlush_valid && LoadQueuePlugin_logic_loadQueue_slots_1_valid) && (((_zz_when_LoadQueuePlugin_l508_4 == _zz_when_LoadQueuePlugin_l508_6) && (_zz_when_LoadQueuePlugin_l508_7 <= _zz_when_LoadQueuePlugin_l508_5)) || ((_zz_when_LoadQueuePlugin_l508_4 != _zz_when_LoadQueuePlugin_l508_6) && (_zz_when_LoadQueuePlugin_l508_5 < _zz_when_LoadQueuePlugin_l508_7))));
  assign _zz_when_LoadQueuePlugin_l508_8 = LoadQueuePlugin_logic_loadQueue_slots_2_robPtr[3];
  assign _zz_when_LoadQueuePlugin_l508_9 = LoadQueuePlugin_logic_loadQueue_slots_2_robPtr[2 : 0];
  assign _zz_when_LoadQueuePlugin_l508_10 = LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr[3];
  assign _zz_when_LoadQueuePlugin_l508_11 = LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr[2 : 0];
  assign when_LoadQueuePlugin_l508_2 = ((LoadQueuePlugin_logic_loadQueue_registeredFlush_valid && LoadQueuePlugin_logic_loadQueue_slots_2_valid) && (((_zz_when_LoadQueuePlugin_l508_8 == _zz_when_LoadQueuePlugin_l508_10) && (_zz_when_LoadQueuePlugin_l508_11 <= _zz_when_LoadQueuePlugin_l508_9)) || ((_zz_when_LoadQueuePlugin_l508_8 != _zz_when_LoadQueuePlugin_l508_10) && (_zz_when_LoadQueuePlugin_l508_9 < _zz_when_LoadQueuePlugin_l508_11))));
  assign _zz_when_LoadQueuePlugin_l508_12 = LoadQueuePlugin_logic_loadQueue_slots_3_robPtr[3];
  assign _zz_when_LoadQueuePlugin_l508_13 = LoadQueuePlugin_logic_loadQueue_slots_3_robPtr[2 : 0];
  assign _zz_when_LoadQueuePlugin_l508_14 = LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr[3];
  assign _zz_when_LoadQueuePlugin_l508_15 = LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr[2 : 0];
  assign when_LoadQueuePlugin_l508_3 = ((LoadQueuePlugin_logic_loadQueue_registeredFlush_valid && LoadQueuePlugin_logic_loadQueue_slots_3_valid) && (((_zz_when_LoadQueuePlugin_l508_12 == _zz_when_LoadQueuePlugin_l508_14) && (_zz_when_LoadQueuePlugin_l508_15 <= _zz_when_LoadQueuePlugin_l508_13)) || ((_zz_when_LoadQueuePlugin_l508_12 != _zz_when_LoadQueuePlugin_l508_14) && (_zz_when_LoadQueuePlugin_l508_13 < _zz_when_LoadQueuePlugin_l508_15))));
  assign AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp = ((AluIntEU_AluIntEuPlugin_gprReadPorts_0_address == 6'h0) ? 32'h0 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp);
  assign AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp = ((AluIntEU_AluIntEuPlugin_gprReadPorts_1_address == 6'h0) ? 32'h0 : _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp);
  assign MulEU_MulEuPlugin_gprReadPorts_0_rsp = ((MulEU_MulEuPlugin_gprReadPorts_0_address == 6'h0) ? 32'h0 : _zz_MulEU_MulEuPlugin_gprReadPorts_0_rsp);
  assign MulEU_MulEuPlugin_gprReadPorts_1_rsp = ((MulEU_MulEuPlugin_gprReadPorts_1_address == 6'h0) ? 32'h0 : _zz_MulEU_MulEuPlugin_gprReadPorts_1_rsp);
  assign BranchEU_BranchEuPlugin_gprReadPorts_0_rsp = ((BranchEU_BranchEuPlugin_gprReadPorts_0_address == 6'h0) ? 32'h0 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_rsp);
  assign BranchEU_BranchEuPlugin_gprReadPorts_1_rsp = ((BranchEU_BranchEuPlugin_gprReadPorts_1_address == 6'h0) ? 32'h0 : _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_rsp);
  assign LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp = ((LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_address == 6'h0) ? 32'h0 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp);
  assign LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp = ((LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_address == 6'h0) ? 32'h0 : _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp);
  assign when_PhysicalRegFile_l130 = (AluIntEU_AluIntEuPlugin_gprWritePort_valid && (AluIntEU_AluIntEuPlugin_gprWritePort_address != 6'h0));
  assign _zz_58 = ({63'd0,1'b1} <<< AluIntEU_AluIntEuPlugin_gprWritePort_address);
  assign when_PhysicalRegFile_l130_1 = (MulEU_MulEuPlugin_gprWritePort_valid && (MulEU_MulEuPlugin_gprWritePort_address != 6'h0));
  assign _zz_59 = ({63'd0,1'b1} <<< MulEU_MulEuPlugin_gprWritePort_address);
  assign when_PhysicalRegFile_l130_2 = (BranchEU_BranchEuPlugin_gprWritePort_valid && (BranchEU_BranchEuPlugin_gprWritePort_address != 6'h0));
  assign _zz_60 = ({63'd0,1'b1} <<< BranchEU_BranchEuPlugin_gprWritePort_address);
  assign when_PhysicalRegFile_l130_3 = (LsuEU_LsuEuPlugin_gprWritePort_valid && (LsuEU_LsuEuPlugin_gprWritePort_address != 6'h0));
  assign _zz_61 = ({63'd0,1'b1} <<< LsuEU_LsuEuPlugin_gprWritePort_address);
  assign when_PhysicalRegFile_l130_4 = (LoadQueuePlugin_hw_prfWritePort_valid && (LoadQueuePlugin_hw_prfWritePort_address != 6'h0));
  assign _zz_62 = ({63'd0,1'b1} <<< LoadQueuePlugin_hw_prfWritePort_address);
  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush = StoreBufferPlugin_logic_slots_0_isFlush;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_addr = StoreBufferPlugin_logic_slots_0_addr;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_addr = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_addr;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_addr = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_data = StoreBufferPlugin_logic_slots_0_data;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_data = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_data;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_data = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_be = StoreBufferPlugin_logic_slots_0_be;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_be = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_be;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_be = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr = StoreBufferPlugin_logic_slots_0_robPtr;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize = StoreBufferPlugin_logic_slots_0_accessSize;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize = MemAccessSize_W;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO = StoreBufferPlugin_logic_slots_0_isIO;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_valid = StoreBufferPlugin_logic_slots_0_valid;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_valid = 1'b1;
      end
    end
    if(when_StoreBufferPlugin_l525) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_valid = 1'b0;
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_valid = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException = StoreBufferPlugin_logic_slots_0_hasEarlyException;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException;
      end
    end
    if(StoreBufferPlugin_logic_mmioResponseForHead) begin
      if(CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_payload_error) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException = 1'b1;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode = StoreBufferPlugin_logic_slots_0_earlyExceptionCode;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode;
      end
    end
    if(StoreBufferPlugin_logic_mmioResponseForHead) begin
      if(CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_payload_error) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode = 8'h07;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_isCommitted = StoreBufferPlugin_logic_slots_0_isCommitted;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_isCommitted = 1'b0;
      end
    end
    if(!when_StoreBufferPlugin_l525) begin
      if(when_StoreBufferPlugin_l529) begin
        if(when_StoreBufferPlugin_l533) begin
          StoreBufferPlugin_logic_slotsAfterUpdates_0_isCommitted = 1'b1;
        end
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_isCommitted = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd = StoreBufferPlugin_logic_slots_0_sentCmd;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd = 1'b0;
      end
    end
    if(StoreBufferPlugin_logic_dcacheCmdFired) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd = 1'b1;
    end
    if(StoreBufferPlugin_logic_mmioCmdFired) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd = 1'b1;
    end
    if(StoreBufferPlugin_logic_dcacheResponseForHead) begin
      if(StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_redo) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd = 1'b0;
      end
    end
    if(StoreBufferPlugin_logic_waitedRefillIsDone) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd = 1'b0;
    end
    if(when_StoreBufferPlugin_l474) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd = 1'b0;
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp = StoreBufferPlugin_logic_slots_0_waitRsp;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp = 1'b0;
      end
    end
    if(StoreBufferPlugin_logic_dcacheCmdFired) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp = 1'b1;
    end
    if(StoreBufferPlugin_logic_mmioCmdFired) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp = 1'b1;
    end
    if(StoreBufferPlugin_logic_dcacheResponseForHead) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp = 1'b0;
    end
    if(StoreBufferPlugin_logic_mmioResponseForHead) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp = 1'b0;
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForRefill = StoreBufferPlugin_logic_slots_0_isWaitingForRefill;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForRefill = 1'b0;
      end
    end
    if(StoreBufferPlugin_logic_dcacheResponseForHead) begin
      if(StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_redo) begin
        if(!StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_flush) begin
          StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForRefill = 1'b1;
        end
      end
    end
    if(StoreBufferPlugin_logic_waitedRefillIsDone) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForRefill = 1'b0;
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForRefill = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForWb = StoreBufferPlugin_logic_slots_0_isWaitingForWb;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForWb = 1'b0;
      end
    end
    if(StoreBufferPlugin_logic_dcacheResponseForHead) begin
      if(StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_redo) begin
        if(StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_flush) begin
          StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForWb = 1'b1;
        end
      end
    end
    if(when_StoreBufferPlugin_l474) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForWb = 1'b0;
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForWb = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_0_refillSlotToWatch = StoreBufferPlugin_logic_slots_0_refillSlotToWatch;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_66) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_0_refillSlotToWatch = 8'h0;
      end
    end
    if(StoreBufferPlugin_logic_dcacheResponseForHead) begin
      if(StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_redo) begin
        if(!StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_flush) begin
          StoreBufferPlugin_logic_slotsAfterUpdates_0_refillSlotToWatch = StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_refillSlot;
        end
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_0_refillSlotToWatch = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_isFlush = StoreBufferPlugin_logic_slots_1_isFlush;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_isFlush = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_isFlush = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_addr = StoreBufferPlugin_logic_slots_1_addr;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_addr = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_addr;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_addr = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_data = StoreBufferPlugin_logic_slots_1_data;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_data = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_data;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_data = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_be = StoreBufferPlugin_logic_slots_1_be;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_be = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_be;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_be = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_robPtr = StoreBufferPlugin_logic_slots_1_robPtr;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_robPtr = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize = StoreBufferPlugin_logic_slots_1_accessSize;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize = MemAccessSize_W;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_isIO = StoreBufferPlugin_logic_slots_1_isIO;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_isIO = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_isIO = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_valid = StoreBufferPlugin_logic_slots_1_valid;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_valid = 1'b1;
      end
    end
    if(when_StoreBufferPlugin_l525_1) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_valid = 1'b0;
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_valid = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_hasEarlyException = StoreBufferPlugin_logic_slots_1_hasEarlyException;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_hasEarlyException = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_hasEarlyException = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_earlyExceptionCode = StoreBufferPlugin_logic_slots_1_earlyExceptionCode;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_earlyExceptionCode = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_earlyExceptionCode = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_isCommitted = StoreBufferPlugin_logic_slots_1_isCommitted;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_isCommitted = 1'b0;
      end
    end
    if(!when_StoreBufferPlugin_l525_1) begin
      if(when_StoreBufferPlugin_l529_1) begin
        if(when_StoreBufferPlugin_l533_1) begin
          StoreBufferPlugin_logic_slotsAfterUpdates_1_isCommitted = 1'b1;
        end
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_isCommitted = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_sentCmd = StoreBufferPlugin_logic_slots_1_sentCmd;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_sentCmd = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_sentCmd = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_waitRsp = StoreBufferPlugin_logic_slots_1_waitRsp;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_waitRsp = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_waitRsp = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForRefill = StoreBufferPlugin_logic_slots_1_isWaitingForRefill;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForRefill = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForRefill = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForWb = StoreBufferPlugin_logic_slots_1_isWaitingForWb;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForWb = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForWb = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_1_refillSlotToWatch = StoreBufferPlugin_logic_slots_1_refillSlotToWatch;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_67) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_1_refillSlotToWatch = 8'h0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_1_refillSlotToWatch = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_isFlush = StoreBufferPlugin_logic_slots_2_isFlush;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_isFlush = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_isFlush = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_addr = StoreBufferPlugin_logic_slots_2_addr;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_addr = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_addr;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_addr = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_data = StoreBufferPlugin_logic_slots_2_data;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_data = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_data;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_data = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_be = StoreBufferPlugin_logic_slots_2_be;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_be = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_be;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_be = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_robPtr = StoreBufferPlugin_logic_slots_2_robPtr;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_robPtr = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize = StoreBufferPlugin_logic_slots_2_accessSize;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize = MemAccessSize_W;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_isIO = StoreBufferPlugin_logic_slots_2_isIO;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_isIO = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_isIO = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_valid = StoreBufferPlugin_logic_slots_2_valid;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_valid = 1'b1;
      end
    end
    if(when_StoreBufferPlugin_l525_2) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_valid = 1'b0;
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_valid = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_hasEarlyException = StoreBufferPlugin_logic_slots_2_hasEarlyException;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_hasEarlyException = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_hasEarlyException = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_earlyExceptionCode = StoreBufferPlugin_logic_slots_2_earlyExceptionCode;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_earlyExceptionCode = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_earlyExceptionCode = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_isCommitted = StoreBufferPlugin_logic_slots_2_isCommitted;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_isCommitted = 1'b0;
      end
    end
    if(!when_StoreBufferPlugin_l525_2) begin
      if(when_StoreBufferPlugin_l529_2) begin
        if(when_StoreBufferPlugin_l533_2) begin
          StoreBufferPlugin_logic_slotsAfterUpdates_2_isCommitted = 1'b1;
        end
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_isCommitted = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_sentCmd = StoreBufferPlugin_logic_slots_2_sentCmd;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_sentCmd = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_sentCmd = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_waitRsp = StoreBufferPlugin_logic_slots_2_waitRsp;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_waitRsp = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_waitRsp = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForRefill = StoreBufferPlugin_logic_slots_2_isWaitingForRefill;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForRefill = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForRefill = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForWb = StoreBufferPlugin_logic_slots_2_isWaitingForWb;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForWb = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForWb = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_2_refillSlotToWatch = StoreBufferPlugin_logic_slots_2_refillSlotToWatch;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_68) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_2_refillSlotToWatch = 8'h0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_2_refillSlotToWatch = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_isFlush = StoreBufferPlugin_logic_slots_3_isFlush;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_isFlush = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_isFlush = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_addr = StoreBufferPlugin_logic_slots_3_addr;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_addr = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_addr;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_addr = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_data = StoreBufferPlugin_logic_slots_3_data;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_data = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_data;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_data = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_be = StoreBufferPlugin_logic_slots_3_be;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_be = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_be;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_be = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_robPtr = StoreBufferPlugin_logic_slots_3_robPtr;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_robPtr = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize = StoreBufferPlugin_logic_slots_3_accessSize;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize = MemAccessSize_W;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_isIO = StoreBufferPlugin_logic_slots_3_isIO;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_isIO = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_isIO = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_valid = StoreBufferPlugin_logic_slots_3_valid;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_valid = 1'b1;
      end
    end
    if(when_StoreBufferPlugin_l525_3) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_valid = 1'b0;
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_valid = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_hasEarlyException = StoreBufferPlugin_logic_slots_3_hasEarlyException;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_hasEarlyException = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_hasEarlyException = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_earlyExceptionCode = StoreBufferPlugin_logic_slots_3_earlyExceptionCode;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_earlyExceptionCode = _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_earlyExceptionCode = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_isCommitted = StoreBufferPlugin_logic_slots_3_isCommitted;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_isCommitted = 1'b0;
      end
    end
    if(!when_StoreBufferPlugin_l525_3) begin
      if(when_StoreBufferPlugin_l529_3) begin
        if(when_StoreBufferPlugin_l533_3) begin
          StoreBufferPlugin_logic_slotsAfterUpdates_3_isCommitted = 1'b1;
        end
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_isCommitted = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_sentCmd = StoreBufferPlugin_logic_slots_3_sentCmd;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_sentCmd = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_sentCmd = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_waitRsp = StoreBufferPlugin_logic_slots_3_waitRsp;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_waitRsp = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_waitRsp = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForRefill = StoreBufferPlugin_logic_slots_3_isWaitingForRefill;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForRefill = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForRefill = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForWb = StoreBufferPlugin_logic_slots_3_isWaitingForWb;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForWb = 1'b0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForWb = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsAfterUpdates_3_refillSlotToWatch = StoreBufferPlugin_logic_slots_3_refillSlotToWatch;
    if(StoreBufferPlugin_hw_pushPortInst_fire) begin
      if(_zz_69) begin
        StoreBufferPlugin_logic_slotsAfterUpdates_3_refillSlotToWatch = 8'h0;
      end
    end
    if(when_StoreBufferPlugin_l540) begin
      StoreBufferPlugin_logic_slotsAfterUpdates_3_refillSlotToWatch = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_isFlush = StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_isFlush = StoreBufferPlugin_logic_slotsAfterUpdates_1_isFlush;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_addr = StoreBufferPlugin_logic_slotsAfterUpdates_0_addr;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_addr = StoreBufferPlugin_logic_slotsAfterUpdates_1_addr;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_data = StoreBufferPlugin_logic_slotsAfterUpdates_0_data;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_data = StoreBufferPlugin_logic_slotsAfterUpdates_1_data;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_be = StoreBufferPlugin_logic_slotsAfterUpdates_0_be;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_be = StoreBufferPlugin_logic_slotsAfterUpdates_1_be;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_robPtr = StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_robPtr = StoreBufferPlugin_logic_slotsAfterUpdates_1_robPtr;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_accessSize = StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_accessSize = StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_isIO = StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_isIO = StoreBufferPlugin_logic_slotsAfterUpdates_1_isIO;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_valid = StoreBufferPlugin_logic_slotsAfterUpdates_0_valid;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_valid = StoreBufferPlugin_logic_slotsAfterUpdates_1_valid;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_hasEarlyException = StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_hasEarlyException = StoreBufferPlugin_logic_slotsAfterUpdates_1_hasEarlyException;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_earlyExceptionCode = StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_earlyExceptionCode = StoreBufferPlugin_logic_slotsAfterUpdates_1_earlyExceptionCode;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_isCommitted = StoreBufferPlugin_logic_slotsAfterUpdates_0_isCommitted;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_isCommitted = StoreBufferPlugin_logic_slotsAfterUpdates_1_isCommitted;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_sentCmd = StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_sentCmd = StoreBufferPlugin_logic_slotsAfterUpdates_1_sentCmd;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_waitRsp = StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_waitRsp = StoreBufferPlugin_logic_slotsAfterUpdates_1_waitRsp;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_isWaitingForRefill = StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForRefill;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_isWaitingForRefill = StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForRefill;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_isWaitingForWb = StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForWb;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_isWaitingForWb = StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForWb;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_0_refillSlotToWatch = StoreBufferPlugin_logic_slotsAfterUpdates_0_refillSlotToWatch;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_0_refillSlotToWatch = StoreBufferPlugin_logic_slotsAfterUpdates_1_refillSlotToWatch;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_isFlush = StoreBufferPlugin_logic_slotsAfterUpdates_1_isFlush;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_isFlush = StoreBufferPlugin_logic_slotsAfterUpdates_2_isFlush;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_addr = StoreBufferPlugin_logic_slotsAfterUpdates_1_addr;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_addr = StoreBufferPlugin_logic_slotsAfterUpdates_2_addr;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_data = StoreBufferPlugin_logic_slotsAfterUpdates_1_data;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_data = StoreBufferPlugin_logic_slotsAfterUpdates_2_data;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_be = StoreBufferPlugin_logic_slotsAfterUpdates_1_be;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_be = StoreBufferPlugin_logic_slotsAfterUpdates_2_be;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_robPtr = StoreBufferPlugin_logic_slotsAfterUpdates_1_robPtr;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_robPtr = StoreBufferPlugin_logic_slotsAfterUpdates_2_robPtr;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_accessSize = StoreBufferPlugin_logic_slotsAfterUpdates_1_accessSize;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_accessSize = StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_isIO = StoreBufferPlugin_logic_slotsAfterUpdates_1_isIO;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_isIO = StoreBufferPlugin_logic_slotsAfterUpdates_2_isIO;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_valid = StoreBufferPlugin_logic_slotsAfterUpdates_1_valid;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_valid = StoreBufferPlugin_logic_slotsAfterUpdates_2_valid;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_hasEarlyException = StoreBufferPlugin_logic_slotsAfterUpdates_1_hasEarlyException;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_hasEarlyException = StoreBufferPlugin_logic_slotsAfterUpdates_2_hasEarlyException;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_earlyExceptionCode = StoreBufferPlugin_logic_slotsAfterUpdates_1_earlyExceptionCode;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_earlyExceptionCode = StoreBufferPlugin_logic_slotsAfterUpdates_2_earlyExceptionCode;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_isCommitted = StoreBufferPlugin_logic_slotsAfterUpdates_1_isCommitted;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_isCommitted = StoreBufferPlugin_logic_slotsAfterUpdates_2_isCommitted;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_sentCmd = StoreBufferPlugin_logic_slotsAfterUpdates_1_sentCmd;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_sentCmd = StoreBufferPlugin_logic_slotsAfterUpdates_2_sentCmd;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_waitRsp = StoreBufferPlugin_logic_slotsAfterUpdates_1_waitRsp;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_waitRsp = StoreBufferPlugin_logic_slotsAfterUpdates_2_waitRsp;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_isWaitingForRefill = StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForRefill;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_isWaitingForRefill = StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForRefill;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_isWaitingForWb = StoreBufferPlugin_logic_slotsAfterUpdates_1_isWaitingForWb;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_isWaitingForWb = StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForWb;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_1_refillSlotToWatch = StoreBufferPlugin_logic_slotsAfterUpdates_1_refillSlotToWatch;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_1_refillSlotToWatch = StoreBufferPlugin_logic_slotsAfterUpdates_2_refillSlotToWatch;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_isFlush = StoreBufferPlugin_logic_slotsAfterUpdates_2_isFlush;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_isFlush = StoreBufferPlugin_logic_slotsAfterUpdates_3_isFlush;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_addr = StoreBufferPlugin_logic_slotsAfterUpdates_2_addr;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_addr = StoreBufferPlugin_logic_slotsAfterUpdates_3_addr;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_data = StoreBufferPlugin_logic_slotsAfterUpdates_2_data;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_data = StoreBufferPlugin_logic_slotsAfterUpdates_3_data;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_be = StoreBufferPlugin_logic_slotsAfterUpdates_2_be;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_be = StoreBufferPlugin_logic_slotsAfterUpdates_3_be;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_robPtr = StoreBufferPlugin_logic_slotsAfterUpdates_2_robPtr;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_robPtr = StoreBufferPlugin_logic_slotsAfterUpdates_3_robPtr;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_accessSize = StoreBufferPlugin_logic_slotsAfterUpdates_2_accessSize;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_accessSize = StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_isIO = StoreBufferPlugin_logic_slotsAfterUpdates_2_isIO;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_isIO = StoreBufferPlugin_logic_slotsAfterUpdates_3_isIO;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_valid = StoreBufferPlugin_logic_slotsAfterUpdates_2_valid;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_valid = StoreBufferPlugin_logic_slotsAfterUpdates_3_valid;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_hasEarlyException = StoreBufferPlugin_logic_slotsAfterUpdates_2_hasEarlyException;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_hasEarlyException = StoreBufferPlugin_logic_slotsAfterUpdates_3_hasEarlyException;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_earlyExceptionCode = StoreBufferPlugin_logic_slotsAfterUpdates_2_earlyExceptionCode;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_earlyExceptionCode = StoreBufferPlugin_logic_slotsAfterUpdates_3_earlyExceptionCode;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_isCommitted = StoreBufferPlugin_logic_slotsAfterUpdates_2_isCommitted;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_isCommitted = StoreBufferPlugin_logic_slotsAfterUpdates_3_isCommitted;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_sentCmd = StoreBufferPlugin_logic_slotsAfterUpdates_2_sentCmd;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_sentCmd = StoreBufferPlugin_logic_slotsAfterUpdates_3_sentCmd;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_waitRsp = StoreBufferPlugin_logic_slotsAfterUpdates_2_waitRsp;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_waitRsp = StoreBufferPlugin_logic_slotsAfterUpdates_3_waitRsp;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_isWaitingForRefill = StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForRefill;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_isWaitingForRefill = StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForRefill;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_isWaitingForWb = StoreBufferPlugin_logic_slotsAfterUpdates_2_isWaitingForWb;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_isWaitingForWb = StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForWb;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_2_refillSlotToWatch = StoreBufferPlugin_logic_slotsAfterUpdates_2_refillSlotToWatch;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_2_refillSlotToWatch = StoreBufferPlugin_logic_slotsAfterUpdates_3_refillSlotToWatch;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_isFlush = StoreBufferPlugin_logic_slotsAfterUpdates_3_isFlush;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_isFlush = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_addr = StoreBufferPlugin_logic_slotsAfterUpdates_3_addr;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_addr = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_data = StoreBufferPlugin_logic_slotsAfterUpdates_3_data;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_data = 32'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_be = StoreBufferPlugin_logic_slotsAfterUpdates_3_be;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_be = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_robPtr = StoreBufferPlugin_logic_slotsAfterUpdates_3_robPtr;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_robPtr = 4'b0000;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_accessSize = StoreBufferPlugin_logic_slotsAfterUpdates_3_accessSize;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_accessSize = MemAccessSize_W;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_isIO = StoreBufferPlugin_logic_slotsAfterUpdates_3_isIO;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_isIO = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_valid = StoreBufferPlugin_logic_slotsAfterUpdates_3_valid;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_valid = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_hasEarlyException = StoreBufferPlugin_logic_slotsAfterUpdates_3_hasEarlyException;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_hasEarlyException = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_earlyExceptionCode = StoreBufferPlugin_logic_slotsAfterUpdates_3_earlyExceptionCode;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_earlyExceptionCode = 8'h0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_isCommitted = StoreBufferPlugin_logic_slotsAfterUpdates_3_isCommitted;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_isCommitted = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_sentCmd = StoreBufferPlugin_logic_slotsAfterUpdates_3_sentCmd;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_sentCmd = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_waitRsp = StoreBufferPlugin_logic_slotsAfterUpdates_3_waitRsp;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_waitRsp = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_isWaitingForRefill = StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForRefill;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_isWaitingForRefill = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_isWaitingForWb = StoreBufferPlugin_logic_slotsAfterUpdates_3_isWaitingForWb;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_isWaitingForWb = 1'b0;
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_slotsNext_3_refillSlotToWatch = StoreBufferPlugin_logic_slotsAfterUpdates_3_refillSlotToWatch;
    if(StoreBufferPlugin_logic_popRequest) begin
      StoreBufferPlugin_logic_slotsNext_3_refillSlotToWatch = 8'h0;
    end
  end

  assign StoreBufferPlugin_logic_flushInProgress = (ROBPlugin_aggregatedFlushSignal_valid && (ROBPlugin_aggregatedFlushSignal_payload_reason == FlushReason_ROLLBACK_TO_ROB_IDX));
  assign StoreBufferPlugin_logic_validFall_0 = (! StoreBufferPlugin_logic_slots_0_valid);
  assign StoreBufferPlugin_logic_validFall_1 = (StoreBufferPlugin_logic_slots_0_valid && (! StoreBufferPlugin_logic_slots_1_valid));
  assign StoreBufferPlugin_logic_validFall_2 = (StoreBufferPlugin_logic_slots_1_valid && (! StoreBufferPlugin_logic_slots_2_valid));
  assign StoreBufferPlugin_logic_validFall_3 = (StoreBufferPlugin_logic_slots_2_valid && (! StoreBufferPlugin_logic_slots_3_valid));
  assign StoreBufferPlugin_logic_canPush = ((|{StoreBufferPlugin_logic_validFall_3,{StoreBufferPlugin_logic_validFall_2,{StoreBufferPlugin_logic_validFall_1,StoreBufferPlugin_logic_validFall_0}}}) && (! StoreBufferPlugin_logic_flushInProgress));
  assign StoreBufferPlugin_hw_pushPortInst_ready = StoreBufferPlugin_logic_canPush;
  assign _zz_63 = (StoreBufferPlugin_logic_validFall_1 || StoreBufferPlugin_logic_validFall_3);
  assign _zz_64 = (StoreBufferPlugin_logic_validFall_2 || StoreBufferPlugin_logic_validFall_3);
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush = StoreBufferPlugin_hw_pushPortInst_payload_isFlush;
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_addr = StoreBufferPlugin_hw_pushPortInst_payload_addr;
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_data = StoreBufferPlugin_hw_pushPortInst_payload_data;
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_be = StoreBufferPlugin_hw_pushPortInst_payload_be;
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr = StoreBufferPlugin_hw_pushPortInst_payload_robPtr;
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_accessSize = StoreBufferPlugin_hw_pushPortInst_payload_accessSize;
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO = StoreBufferPlugin_hw_pushPortInst_payload_isIO;
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException = StoreBufferPlugin_hw_pushPortInst_payload_hasEarlyException;
  assign _zz_StoreBufferPlugin_logic_slotsAfterUpdates_0_earlyExceptionCode = StoreBufferPlugin_hw_pushPortInst_payload_earlyExceptionCode;
  assign _zz_65 = ({3'd0,1'b1} <<< {_zz_64,_zz_63});
  assign _zz_66 = _zz_65[0];
  assign _zz_67 = _zz_65[1];
  assign _zz_68 = _zz_65[2];
  assign _zz_69 = _zz_65[3];
  assign StoreBufferPlugin_logic_sharedWriteCond = ((((((StoreBufferPlugin_logic_slots_0_valid && StoreBufferPlugin_logic_slots_0_isCommitted) && (! StoreBufferPlugin_logic_slots_0_isFlush)) && (! StoreBufferPlugin_logic_slots_0_waitRsp)) && (! StoreBufferPlugin_logic_slots_0_isWaitingForRefill)) && (! StoreBufferPlugin_logic_slots_0_isWaitingForWb)) && (! StoreBufferPlugin_logic_slots_0_hasEarlyException));
  assign StoreBufferPlugin_logic_canPopNormalOp = (StoreBufferPlugin_logic_sharedWriteCond && (! StoreBufferPlugin_logic_slots_0_isIO));
  assign StoreBufferPlugin_logic_canPopFlushOp = (((StoreBufferPlugin_logic_slots_0_valid && StoreBufferPlugin_logic_slots_0_isFlush) && (! StoreBufferPlugin_logic_slots_0_waitRsp)) && (! StoreBufferPlugin_logic_slots_0_isWaitingForWb));
  assign StoreBufferPlugin_logic_canPopMMIOOp = (StoreBufferPlugin_logic_sharedWriteCond && StoreBufferPlugin_logic_slots_0_isIO);
  assign when_StoreBufferPlugin_l316 = (1'b0 && StoreBufferPlugin_logic_slots_0_isIO);
  assign StoreBufferPlugin_logic_canSendToDCache = (StoreBufferPlugin_logic_canPopNormalOp || StoreBufferPlugin_logic_canPopFlushOp);
  assign StoreBufferPlugin_hw_dCacheStorePort_cmd_valid = StoreBufferPlugin_logic_canSendToDCache;
  always @(*) begin
    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(StoreBufferPlugin_logic_canSendToDCache) begin
      if(StoreBufferPlugin_logic_slots_0_isFlush) begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_address = StoreBufferPlugin_logic_slots_0_addr;
      end else begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_address = StoreBufferPlugin_logic_slots_0_addr;
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(StoreBufferPlugin_logic_canSendToDCache) begin
      if(StoreBufferPlugin_logic_slots_0_isFlush) begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_data = 32'h0;
      end else begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_data = StoreBufferPlugin_logic_slots_0_data;
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_mask = 4'bxxxx;
    if(StoreBufferPlugin_logic_canSendToDCache) begin
      if(StoreBufferPlugin_logic_slots_0_isFlush) begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_mask = 4'b0000;
      end else begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_mask = StoreBufferPlugin_logic_slots_0_be;
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_io = 1'bx;
    if(StoreBufferPlugin_logic_canSendToDCache) begin
      if(StoreBufferPlugin_logic_slots_0_isFlush) begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_io = 1'b0;
      end else begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_io = StoreBufferPlugin_logic_slots_0_isIO;
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flush = 1'bx;
    if(StoreBufferPlugin_logic_canSendToDCache) begin
      if(StoreBufferPlugin_logic_slots_0_isFlush) begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flush = 1'b1;
      end else begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flush = 1'b0;
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flushFree = 1'bx;
    if(StoreBufferPlugin_logic_canSendToDCache) begin
      if(StoreBufferPlugin_logic_slots_0_isFlush) begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flushFree = 1'b0;
      end else begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_flushFree = 1'b0;
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_prefetch = 1'bx;
    if(StoreBufferPlugin_logic_canSendToDCache) begin
      if(StoreBufferPlugin_logic_slots_0_isFlush) begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_prefetch = 1'b0;
      end else begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_prefetch = 1'b0;
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_id = 3'bxxx;
    if(StoreBufferPlugin_logic_canSendToDCache) begin
      if(StoreBufferPlugin_logic_slots_0_isFlush) begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_id = StoreBufferPlugin_logic_slots_0_robPtr[2:0];
      end else begin
        StoreBufferPlugin_hw_dCacheStorePort_cmd_payload_id = StoreBufferPlugin_logic_slots_0_robPtr[2:0];
      end
    end
  end

  assign StoreBufferPlugin_logic_dcacheCmdFired = (StoreBufferPlugin_logic_canSendToDCache && StoreBufferPlugin_hw_dCacheStorePort_cmd_ready);
  assign StoreBufferPlugin_logic_mmioCmdFired = (StoreBufferPlugin_logic_canPopMMIOOp && CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_cmd_ready);
  assign StoreBufferPlugin_logic_dcacheResponseForHead = ((((StoreBufferPlugin_hw_dCacheStorePort_rsp_valid && StoreBufferPlugin_logic_slots_0_valid) && (StoreBufferPlugin_logic_slots_0_waitRsp || StoreBufferPlugin_logic_dcacheCmdFired)) && (! StoreBufferPlugin_logic_slots_0_isIO)) && (_zz_StoreBufferPlugin_logic_dcacheResponseForHead == StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_id));
  assign StoreBufferPlugin_logic_mmioResponseForHead = ((((CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_valid && StoreBufferPlugin_logic_slots_0_valid) && StoreBufferPlugin_logic_slots_0_isIO) && (StoreBufferPlugin_logic_slots_0_waitRsp || StoreBufferPlugin_logic_mmioCmdFired)) && (StoreBufferPlugin_logic_slots_0_robPtr == CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_payload_id));
  assign oneShot_25_io_triggerIn = (StoreBufferPlugin_logic_mmioResponseForHead && (_zz_when_Debug_l71 < _zz_io_triggerIn_22));
  assign _zz_when_Debug_l71_12 = 6'h20;
  assign when_Debug_l71_11 = (_zz_when_Debug_l71 < _zz_when_Debug_l71_11_1);
  assign StoreBufferPlugin_logic_waitedRefillIsDone = ((StoreBufferPlugin_logic_slots_0_valid && StoreBufferPlugin_logic_slots_0_isWaitingForRefill) && (|(StoreBufferPlugin_logic_slots_0_refillSlotToWatch & DataCachePlugin_setup_refillCompletions)));
  assign when_StoreBufferPlugin_l474 = ((StoreBufferPlugin_logic_slots_0_valid && StoreBufferPlugin_logic_slots_0_isWaitingForWb) && (! DataCachePlugin_setup_writebackBusy));
  always @(*) begin
    StoreBufferPlugin_logic_commitUpdateInfo_validMask = 4'b0000;
    StoreBufferPlugin_logic_commitUpdateInfo_validMask[0] = _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask;
    StoreBufferPlugin_logic_commitUpdateInfo_validMask[1] = _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_1;
    StoreBufferPlugin_logic_commitUpdateInfo_validMask[2] = _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_2;
    StoreBufferPlugin_logic_commitUpdateInfo_validMask[3] = _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_3;
  end

  always @(*) begin
    _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask = 1'b0;
    if(when_StoreBufferPlugin_l498) begin
      if(when_StoreBufferPlugin_l504) begin
        _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask = 1'b1;
      end
    end
  end

  assign when_StoreBufferPlugin_l498 = (StoreBufferPlugin_logic_slots_0_valid && (! StoreBufferPlugin_logic_slots_0_isCommitted));
  assign when_StoreBufferPlugin_l504 = (((ROBPlugin_robComponent_io_commit_0_canCommit && (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_robPtr == StoreBufferPlugin_logic_slots_0_robPtr)) && ((ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_uopCode == BaseUopCode_STORE) || 1'b0)) && (! ROBPlugin_robComponent_io_commit_0_entry_status_hasException));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_1 = 1'b0;
    if(when_StoreBufferPlugin_l498_1) begin
      if(when_StoreBufferPlugin_l504_1) begin
        _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_1 = 1'b1;
      end
    end
  end

  assign when_StoreBufferPlugin_l498_1 = (StoreBufferPlugin_logic_slots_1_valid && (! StoreBufferPlugin_logic_slots_1_isCommitted));
  assign when_StoreBufferPlugin_l504_1 = (((ROBPlugin_robComponent_io_commit_0_canCommit && (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_robPtr == StoreBufferPlugin_logic_slots_1_robPtr)) && ((ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_uopCode == BaseUopCode_STORE) || 1'b0)) && (! ROBPlugin_robComponent_io_commit_0_entry_status_hasException));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_2 = 1'b0;
    if(when_StoreBufferPlugin_l498_2) begin
      if(when_StoreBufferPlugin_l504_2) begin
        _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_2 = 1'b1;
      end
    end
  end

  assign when_StoreBufferPlugin_l498_2 = (StoreBufferPlugin_logic_slots_2_valid && (! StoreBufferPlugin_logic_slots_2_isCommitted));
  assign when_StoreBufferPlugin_l504_2 = (((ROBPlugin_robComponent_io_commit_0_canCommit && (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_robPtr == StoreBufferPlugin_logic_slots_2_robPtr)) && ((ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_uopCode == BaseUopCode_STORE) || 1'b0)) && (! ROBPlugin_robComponent_io_commit_0_entry_status_hasException));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_3 = 1'b0;
    if(when_StoreBufferPlugin_l498_3) begin
      if(when_StoreBufferPlugin_l504_3) begin
        _zz_StoreBufferPlugin_logic_commitUpdateInfo_validMask_3 = 1'b1;
      end
    end
  end

  assign when_StoreBufferPlugin_l498_3 = (StoreBufferPlugin_logic_slots_3_valid && (! StoreBufferPlugin_logic_slots_3_isCommitted));
  assign when_StoreBufferPlugin_l504_3 = (((ROBPlugin_robComponent_io_commit_0_canCommit && (ROBPlugin_robComponent_io_commit_0_entry_payload_uop_robPtr == StoreBufferPlugin_logic_slots_3_robPtr)) && ((ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_uopCode == BaseUopCode_STORE) || 1'b0)) && (! ROBPlugin_robComponent_io_commit_0_entry_status_hasException));
  assign _zz_when_StoreBufferPlugin_l525 = StoreBufferPlugin_logic_slots_0_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l525_1 = StoreBufferPlugin_logic_slots_0_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l525_2 = StoreBufferPlugin_logic_registeredFlush_targetRobPtr[3];
  assign _zz_when_StoreBufferPlugin_l525_3 = StoreBufferPlugin_logic_registeredFlush_targetRobPtr[2 : 0];
  assign when_StoreBufferPlugin_l525 = (((StoreBufferPlugin_logic_registeredFlush_valid && StoreBufferPlugin_logic_slots_0_valid) && (! StoreBufferPlugin_logic_slots_0_isCommitted)) && (((_zz_when_StoreBufferPlugin_l525 == _zz_when_StoreBufferPlugin_l525_2) && (_zz_when_StoreBufferPlugin_l525_3 <= _zz_when_StoreBufferPlugin_l525_1)) || ((_zz_when_StoreBufferPlugin_l525 != _zz_when_StoreBufferPlugin_l525_2) && (_zz_when_StoreBufferPlugin_l525_1 < _zz_when_StoreBufferPlugin_l525_3))));
  assign when_StoreBufferPlugin_l533 = StoreBufferPlugin_logic_registeredCommitUpdate_validMask[0];
  assign when_StoreBufferPlugin_l529 = (StoreBufferPlugin_logic_slots_0_valid && (! StoreBufferPlugin_logic_slots_0_isCommitted));
  assign _zz_when_StoreBufferPlugin_l525_4 = StoreBufferPlugin_logic_slots_1_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l525_5 = StoreBufferPlugin_logic_slots_1_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l525_6 = StoreBufferPlugin_logic_registeredFlush_targetRobPtr[3];
  assign _zz_when_StoreBufferPlugin_l525_7 = StoreBufferPlugin_logic_registeredFlush_targetRobPtr[2 : 0];
  assign when_StoreBufferPlugin_l525_1 = (((StoreBufferPlugin_logic_registeredFlush_valid && StoreBufferPlugin_logic_slots_1_valid) && (! StoreBufferPlugin_logic_slots_1_isCommitted)) && (((_zz_when_StoreBufferPlugin_l525_4 == _zz_when_StoreBufferPlugin_l525_6) && (_zz_when_StoreBufferPlugin_l525_7 <= _zz_when_StoreBufferPlugin_l525_5)) || ((_zz_when_StoreBufferPlugin_l525_4 != _zz_when_StoreBufferPlugin_l525_6) && (_zz_when_StoreBufferPlugin_l525_5 < _zz_when_StoreBufferPlugin_l525_7))));
  assign when_StoreBufferPlugin_l533_1 = StoreBufferPlugin_logic_registeredCommitUpdate_validMask[1];
  assign when_StoreBufferPlugin_l529_1 = (StoreBufferPlugin_logic_slots_1_valid && (! StoreBufferPlugin_logic_slots_1_isCommitted));
  assign _zz_when_StoreBufferPlugin_l525_8 = StoreBufferPlugin_logic_slots_2_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l525_9 = StoreBufferPlugin_logic_slots_2_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l525_10 = StoreBufferPlugin_logic_registeredFlush_targetRobPtr[3];
  assign _zz_when_StoreBufferPlugin_l525_11 = StoreBufferPlugin_logic_registeredFlush_targetRobPtr[2 : 0];
  assign when_StoreBufferPlugin_l525_2 = (((StoreBufferPlugin_logic_registeredFlush_valid && StoreBufferPlugin_logic_slots_2_valid) && (! StoreBufferPlugin_logic_slots_2_isCommitted)) && (((_zz_when_StoreBufferPlugin_l525_8 == _zz_when_StoreBufferPlugin_l525_10) && (_zz_when_StoreBufferPlugin_l525_11 <= _zz_when_StoreBufferPlugin_l525_9)) || ((_zz_when_StoreBufferPlugin_l525_8 != _zz_when_StoreBufferPlugin_l525_10) && (_zz_when_StoreBufferPlugin_l525_9 < _zz_when_StoreBufferPlugin_l525_11))));
  assign when_StoreBufferPlugin_l533_2 = StoreBufferPlugin_logic_registeredCommitUpdate_validMask[2];
  assign when_StoreBufferPlugin_l529_2 = (StoreBufferPlugin_logic_slots_2_valid && (! StoreBufferPlugin_logic_slots_2_isCommitted));
  assign _zz_when_StoreBufferPlugin_l525_12 = StoreBufferPlugin_logic_slots_3_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l525_13 = StoreBufferPlugin_logic_slots_3_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l525_14 = StoreBufferPlugin_logic_registeredFlush_targetRobPtr[3];
  assign _zz_when_StoreBufferPlugin_l525_15 = StoreBufferPlugin_logic_registeredFlush_targetRobPtr[2 : 0];
  assign when_StoreBufferPlugin_l525_3 = (((StoreBufferPlugin_logic_registeredFlush_valid && StoreBufferPlugin_logic_slots_3_valid) && (! StoreBufferPlugin_logic_slots_3_isCommitted)) && (((_zz_when_StoreBufferPlugin_l525_12 == _zz_when_StoreBufferPlugin_l525_14) && (_zz_when_StoreBufferPlugin_l525_15 <= _zz_when_StoreBufferPlugin_l525_13)) || ((_zz_when_StoreBufferPlugin_l525_12 != _zz_when_StoreBufferPlugin_l525_14) && (_zz_when_StoreBufferPlugin_l525_13 < _zz_when_StoreBufferPlugin_l525_15))));
  assign when_StoreBufferPlugin_l533_3 = StoreBufferPlugin_logic_registeredCommitUpdate_validMask[3];
  assign when_StoreBufferPlugin_l529_3 = (StoreBufferPlugin_logic_slots_3_valid && (! StoreBufferPlugin_logic_slots_3_isCommitted));
  assign when_StoreBufferPlugin_l540 = (ROBPlugin_aggregatedFlushSignal_valid && (ROBPlugin_aggregatedFlushSignal_payload_reason == FlushReason_FULL_FLUSH));
  assign StoreBufferPlugin_logic_operationDone = (((StoreBufferPlugin_logic_slotsAfterUpdates_0_sentCmd && (! StoreBufferPlugin_logic_slotsAfterUpdates_0_waitRsp)) && (! StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForRefill)) && (! StoreBufferPlugin_logic_slotsAfterUpdates_0_isWaitingForWb));
  always @(*) begin
    StoreBufferPlugin_logic_popRequest = 1'b0;
    if(when_StoreBufferPlugin_l555) begin
      if(StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush) begin
        if(StoreBufferPlugin_logic_operationDone) begin
          StoreBufferPlugin_logic_popRequest = 1'b1;
        end
      end else begin
        if(StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException) begin
          StoreBufferPlugin_logic_popRequest = 1'b1;
        end else begin
          if(StoreBufferPlugin_logic_operationDone) begin
            StoreBufferPlugin_logic_popRequest = 1'b1;
          end
        end
      end
    end else begin
      if(when_StoreBufferPlugin_l576) begin
        StoreBufferPlugin_logic_popRequest = 1'b1;
      end
    end
  end

  assign when_StoreBufferPlugin_l555 = (StoreBufferPlugin_logic_slotsAfterUpdates_0_valid && StoreBufferPlugin_logic_slotsAfterUpdates_0_isCommitted);
  assign when_StoreBufferPlugin_l576 = ((! StoreBufferPlugin_logic_slotsAfterUpdates_0_valid) && (! (|{StoreBufferPlugin_logic_slots_3_valid,{StoreBufferPlugin_logic_slots_2_valid,StoreBufferPlugin_logic_slots_1_valid}})));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask = 4'b0000;
    case(StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size)
      MemAccessSize_B : begin
        _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask = _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask;
      end
      MemAccessSize_H : begin
        _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask = _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_2[3:0];
      end
      MemAccessSize_W : begin
        _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask = _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_5[3:0];
      end
      default : begin
        _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask = 4'b1111;
      end
    endcase
  end

  assign _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_1 = _zz__zz_StoreBufferPlugin_logic_forwardingLogic_loadMask_1[1 : 0];
  assign StoreBufferPlugin_logic_forwardingLogic_loadMask = _zz_StoreBufferPlugin_logic_forwardingLogic_loadMask;
  assign StoreBufferPlugin_logic_forwardingLogic_bypassInitial_data = 32'h0;
  assign StoreBufferPlugin_logic_forwardingLogic_bypassInitial_hitMask = 4'b0000;
  always @(*) begin
    _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data = StoreBufferPlugin_logic_forwardingLogic_bypassInitial_data;
    if(when_StoreBufferPlugin_l631) begin
      if(when_StoreBufferPlugin_l638) begin
        if(when_StoreBufferPlugin_l640) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data[7 : 0] = StoreBufferPlugin_logic_slots_3_data[7 : 0];
        end
        if(when_StoreBufferPlugin_l640_1) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data[15 : 8] = StoreBufferPlugin_logic_slots_3_data[15 : 8];
        end
        if(when_StoreBufferPlugin_l640_2) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data[23 : 16] = StoreBufferPlugin_logic_slots_3_data[23 : 16];
        end
        if(when_StoreBufferPlugin_l640_3) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data[31 : 24] = StoreBufferPlugin_logic_slots_3_data[31 : 24];
        end
      end
    end
  end

  always @(*) begin
    _zz_when_StoreBufferPlugin_l640 = StoreBufferPlugin_logic_forwardingLogic_bypassInitial_hitMask;
    if(when_StoreBufferPlugin_l631) begin
      if(when_StoreBufferPlugin_l638) begin
        if(when_StoreBufferPlugin_l640) begin
          _zz_when_StoreBufferPlugin_l640[0] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_1) begin
          _zz_when_StoreBufferPlugin_l640[1] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_2) begin
          _zz_when_StoreBufferPlugin_l640[2] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_3) begin
          _zz_when_StoreBufferPlugin_l640[3] = 1'b1;
        end
      end
    end
  end

  assign _zz_when_StoreBufferPlugin_l631 = StoreBufferPlugin_logic_slots_3_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l631_1 = StoreBufferPlugin_logic_slots_3_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l631_2 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l631_3 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign when_StoreBufferPlugin_l631 = ((((((StoreBufferPlugin_logic_slots_3_valid && (! StoreBufferPlugin_logic_slots_3_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_3_isFlush)) && (! (((_zz_when_StoreBufferPlugin_l631 == _zz_when_StoreBufferPlugin_l631_2) && (_zz_when_StoreBufferPlugin_l631_3 <= _zz_when_StoreBufferPlugin_l631_1)) || ((_zz_when_StoreBufferPlugin_l631 != _zz_when_StoreBufferPlugin_l631_2) && (_zz_when_StoreBufferPlugin_l631_1 < _zz_when_StoreBufferPlugin_l631_3))))) && (! StoreBufferPlugin_logic_slots_3_waitRsp)) && (! StoreBufferPlugin_logic_slots_3_isWaitingForRefill)) && (! StoreBufferPlugin_logic_slots_3_isWaitingForWb));
  assign _zz_when_StoreBufferPlugin_l638 = StoreBufferPlugin_logic_slots_3_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l638_1 = StoreBufferPlugin_logic_slots_3_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l638_2 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l638_3 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign when_StoreBufferPlugin_l638 = (((! StoreBufferPlugin_logic_slots_3_hasEarlyException) && (! (((_zz_when_StoreBufferPlugin_l638 == _zz_when_StoreBufferPlugin_l638_2) && (_zz_when_StoreBufferPlugin_l638_3 <= _zz_when_StoreBufferPlugin_l638_1)) || ((_zz_when_StoreBufferPlugin_l638 != _zz_when_StoreBufferPlugin_l638_2) && (_zz_when_StoreBufferPlugin_l638_1 < _zz_when_StoreBufferPlugin_l638_3))))) && (StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[31 : 2] == StoreBufferPlugin_logic_slots_3_addr[31 : 2]));
  assign when_StoreBufferPlugin_l640 = ((StoreBufferPlugin_logic_slots_3_be[0] && StoreBufferPlugin_logic_forwardingLogic_loadMask[0]) && (! StoreBufferPlugin_logic_forwardingLogic_bypassInitial_hitMask[0]));
  assign when_StoreBufferPlugin_l640_1 = ((StoreBufferPlugin_logic_slots_3_be[1] && StoreBufferPlugin_logic_forwardingLogic_loadMask[1]) && (! StoreBufferPlugin_logic_forwardingLogic_bypassInitial_hitMask[1]));
  assign when_StoreBufferPlugin_l640_2 = ((StoreBufferPlugin_logic_slots_3_be[2] && StoreBufferPlugin_logic_forwardingLogic_loadMask[2]) && (! StoreBufferPlugin_logic_forwardingLogic_bypassInitial_hitMask[2]));
  assign when_StoreBufferPlugin_l640_3 = ((StoreBufferPlugin_logic_slots_3_be[3] && StoreBufferPlugin_logic_forwardingLogic_loadMask[3]) && (! StoreBufferPlugin_logic_forwardingLogic_bypassInitial_hitMask[3]));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_1 = _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data;
    if(when_StoreBufferPlugin_l631_1) begin
      if(when_StoreBufferPlugin_l638_1) begin
        if(when_StoreBufferPlugin_l640_4) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_1[7 : 0] = StoreBufferPlugin_logic_slots_2_data[7 : 0];
        end
        if(when_StoreBufferPlugin_l640_5) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_1[15 : 8] = StoreBufferPlugin_logic_slots_2_data[15 : 8];
        end
        if(when_StoreBufferPlugin_l640_6) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_1[23 : 16] = StoreBufferPlugin_logic_slots_2_data[23 : 16];
        end
        if(when_StoreBufferPlugin_l640_7) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_1[31 : 24] = StoreBufferPlugin_logic_slots_2_data[31 : 24];
        end
      end
    end
  end

  always @(*) begin
    _zz_when_StoreBufferPlugin_l640_1 = _zz_when_StoreBufferPlugin_l640;
    if(when_StoreBufferPlugin_l631_1) begin
      if(when_StoreBufferPlugin_l638_1) begin
        if(when_StoreBufferPlugin_l640_4) begin
          _zz_when_StoreBufferPlugin_l640_1[0] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_5) begin
          _zz_when_StoreBufferPlugin_l640_1[1] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_6) begin
          _zz_when_StoreBufferPlugin_l640_1[2] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_7) begin
          _zz_when_StoreBufferPlugin_l640_1[3] = 1'b1;
        end
      end
    end
  end

  assign _zz_when_StoreBufferPlugin_l631_4 = StoreBufferPlugin_logic_slots_2_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l631_5 = StoreBufferPlugin_logic_slots_2_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l631_6 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l631_7 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign when_StoreBufferPlugin_l631_1 = ((((((StoreBufferPlugin_logic_slots_2_valid && (! StoreBufferPlugin_logic_slots_2_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_2_isFlush)) && (! (((_zz_when_StoreBufferPlugin_l631_4 == _zz_when_StoreBufferPlugin_l631_6) && (_zz_when_StoreBufferPlugin_l631_7 <= _zz_when_StoreBufferPlugin_l631_5)) || ((_zz_when_StoreBufferPlugin_l631_4 != _zz_when_StoreBufferPlugin_l631_6) && (_zz_when_StoreBufferPlugin_l631_5 < _zz_when_StoreBufferPlugin_l631_7))))) && (! StoreBufferPlugin_logic_slots_2_waitRsp)) && (! StoreBufferPlugin_logic_slots_2_isWaitingForRefill)) && (! StoreBufferPlugin_logic_slots_2_isWaitingForWb));
  assign _zz_when_StoreBufferPlugin_l638_4 = StoreBufferPlugin_logic_slots_2_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l638_5 = StoreBufferPlugin_logic_slots_2_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l638_6 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l638_7 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign when_StoreBufferPlugin_l638_1 = (((! StoreBufferPlugin_logic_slots_2_hasEarlyException) && (! (((_zz_when_StoreBufferPlugin_l638_4 == _zz_when_StoreBufferPlugin_l638_6) && (_zz_when_StoreBufferPlugin_l638_7 <= _zz_when_StoreBufferPlugin_l638_5)) || ((_zz_when_StoreBufferPlugin_l638_4 != _zz_when_StoreBufferPlugin_l638_6) && (_zz_when_StoreBufferPlugin_l638_5 < _zz_when_StoreBufferPlugin_l638_7))))) && (StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[31 : 2] == StoreBufferPlugin_logic_slots_2_addr[31 : 2]));
  assign when_StoreBufferPlugin_l640_4 = ((StoreBufferPlugin_logic_slots_2_be[0] && StoreBufferPlugin_logic_forwardingLogic_loadMask[0]) && (! _zz_when_StoreBufferPlugin_l640[0]));
  assign when_StoreBufferPlugin_l640_5 = ((StoreBufferPlugin_logic_slots_2_be[1] && StoreBufferPlugin_logic_forwardingLogic_loadMask[1]) && (! _zz_when_StoreBufferPlugin_l640[1]));
  assign when_StoreBufferPlugin_l640_6 = ((StoreBufferPlugin_logic_slots_2_be[2] && StoreBufferPlugin_logic_forwardingLogic_loadMask[2]) && (! _zz_when_StoreBufferPlugin_l640[2]));
  assign when_StoreBufferPlugin_l640_7 = ((StoreBufferPlugin_logic_slots_2_be[3] && StoreBufferPlugin_logic_forwardingLogic_loadMask[3]) && (! _zz_when_StoreBufferPlugin_l640[3]));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_2 = _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_1;
    if(when_StoreBufferPlugin_l631_2) begin
      if(when_StoreBufferPlugin_l638_2) begin
        if(when_StoreBufferPlugin_l640_8) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_2[7 : 0] = StoreBufferPlugin_logic_slots_1_data[7 : 0];
        end
        if(when_StoreBufferPlugin_l640_9) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_2[15 : 8] = StoreBufferPlugin_logic_slots_1_data[15 : 8];
        end
        if(when_StoreBufferPlugin_l640_10) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_2[23 : 16] = StoreBufferPlugin_logic_slots_1_data[23 : 16];
        end
        if(when_StoreBufferPlugin_l640_11) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_2[31 : 24] = StoreBufferPlugin_logic_slots_1_data[31 : 24];
        end
      end
    end
  end

  always @(*) begin
    _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask = _zz_when_StoreBufferPlugin_l640_1;
    if(when_StoreBufferPlugin_l631_2) begin
      if(when_StoreBufferPlugin_l638_2) begin
        if(when_StoreBufferPlugin_l640_8) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[0] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_9) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[1] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_10) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[2] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_11) begin
          _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[3] = 1'b1;
        end
      end
    end
  end

  assign _zz_when_StoreBufferPlugin_l631_8 = StoreBufferPlugin_logic_slots_1_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l631_9 = StoreBufferPlugin_logic_slots_1_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l631_10 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l631_11 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign when_StoreBufferPlugin_l631_2 = ((((((StoreBufferPlugin_logic_slots_1_valid && (! StoreBufferPlugin_logic_slots_1_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_1_isFlush)) && (! (((_zz_when_StoreBufferPlugin_l631_8 == _zz_when_StoreBufferPlugin_l631_10) && (_zz_when_StoreBufferPlugin_l631_11 <= _zz_when_StoreBufferPlugin_l631_9)) || ((_zz_when_StoreBufferPlugin_l631_8 != _zz_when_StoreBufferPlugin_l631_10) && (_zz_when_StoreBufferPlugin_l631_9 < _zz_when_StoreBufferPlugin_l631_11))))) && (! StoreBufferPlugin_logic_slots_1_waitRsp)) && (! StoreBufferPlugin_logic_slots_1_isWaitingForRefill)) && (! StoreBufferPlugin_logic_slots_1_isWaitingForWb));
  assign _zz_when_StoreBufferPlugin_l638_8 = StoreBufferPlugin_logic_slots_1_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l638_9 = StoreBufferPlugin_logic_slots_1_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l638_10 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l638_11 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign when_StoreBufferPlugin_l638_2 = (((! StoreBufferPlugin_logic_slots_1_hasEarlyException) && (! (((_zz_when_StoreBufferPlugin_l638_8 == _zz_when_StoreBufferPlugin_l638_10) && (_zz_when_StoreBufferPlugin_l638_11 <= _zz_when_StoreBufferPlugin_l638_9)) || ((_zz_when_StoreBufferPlugin_l638_8 != _zz_when_StoreBufferPlugin_l638_10) && (_zz_when_StoreBufferPlugin_l638_9 < _zz_when_StoreBufferPlugin_l638_11))))) && (StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[31 : 2] == StoreBufferPlugin_logic_slots_1_addr[31 : 2]));
  assign when_StoreBufferPlugin_l640_8 = ((StoreBufferPlugin_logic_slots_1_be[0] && StoreBufferPlugin_logic_forwardingLogic_loadMask[0]) && (! _zz_when_StoreBufferPlugin_l640_1[0]));
  assign when_StoreBufferPlugin_l640_9 = ((StoreBufferPlugin_logic_slots_1_be[1] && StoreBufferPlugin_logic_forwardingLogic_loadMask[1]) && (! _zz_when_StoreBufferPlugin_l640_1[1]));
  assign when_StoreBufferPlugin_l640_10 = ((StoreBufferPlugin_logic_slots_1_be[2] && StoreBufferPlugin_logic_forwardingLogic_loadMask[2]) && (! _zz_when_StoreBufferPlugin_l640_1[2]));
  assign when_StoreBufferPlugin_l640_11 = ((StoreBufferPlugin_logic_slots_1_be[3] && StoreBufferPlugin_logic_forwardingLogic_loadMask[3]) && (! _zz_when_StoreBufferPlugin_l640_1[3]));
  always @(*) begin
    StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data = _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data_2;
    if(when_StoreBufferPlugin_l631_3) begin
      if(when_StoreBufferPlugin_l638_3) begin
        if(when_StoreBufferPlugin_l640_12) begin
          StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data[7 : 0] = StoreBufferPlugin_logic_slots_0_data[7 : 0];
        end
        if(when_StoreBufferPlugin_l640_13) begin
          StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data[15 : 8] = StoreBufferPlugin_logic_slots_0_data[15 : 8];
        end
        if(when_StoreBufferPlugin_l640_14) begin
          StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data[23 : 16] = StoreBufferPlugin_logic_slots_0_data[23 : 16];
        end
        if(when_StoreBufferPlugin_l640_15) begin
          StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data[31 : 24] = StoreBufferPlugin_logic_slots_0_data[31 : 24];
        end
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask = _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask;
    if(when_StoreBufferPlugin_l631_3) begin
      if(when_StoreBufferPlugin_l638_3) begin
        if(when_StoreBufferPlugin_l640_12) begin
          StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[0] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_13) begin
          StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[1] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_14) begin
          StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[2] = 1'b1;
        end
        if(when_StoreBufferPlugin_l640_15) begin
          StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[3] = 1'b1;
        end
      end
    end
  end

  assign _zz_when_StoreBufferPlugin_l631_12 = StoreBufferPlugin_logic_slots_0_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l631_13 = StoreBufferPlugin_logic_slots_0_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l631_14 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l631_15 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign when_StoreBufferPlugin_l631_3 = ((((((StoreBufferPlugin_logic_slots_0_valid && (! StoreBufferPlugin_logic_slots_0_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_0_isFlush)) && (! (((_zz_when_StoreBufferPlugin_l631_12 == _zz_when_StoreBufferPlugin_l631_14) && (_zz_when_StoreBufferPlugin_l631_15 <= _zz_when_StoreBufferPlugin_l631_13)) || ((_zz_when_StoreBufferPlugin_l631_12 != _zz_when_StoreBufferPlugin_l631_14) && (_zz_when_StoreBufferPlugin_l631_13 < _zz_when_StoreBufferPlugin_l631_15))))) && (! StoreBufferPlugin_logic_slots_0_waitRsp)) && (! StoreBufferPlugin_logic_slots_0_isWaitingForRefill)) && (! StoreBufferPlugin_logic_slots_0_isWaitingForWb));
  assign _zz_when_StoreBufferPlugin_l638_12 = StoreBufferPlugin_logic_slots_0_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l638_13 = StoreBufferPlugin_logic_slots_0_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l638_14 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l638_15 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign when_StoreBufferPlugin_l638_3 = (((! StoreBufferPlugin_logic_slots_0_hasEarlyException) && (! (((_zz_when_StoreBufferPlugin_l638_12 == _zz_when_StoreBufferPlugin_l638_14) && (_zz_when_StoreBufferPlugin_l638_15 <= _zz_when_StoreBufferPlugin_l638_13)) || ((_zz_when_StoreBufferPlugin_l638_12 != _zz_when_StoreBufferPlugin_l638_14) && (_zz_when_StoreBufferPlugin_l638_13 < _zz_when_StoreBufferPlugin_l638_15))))) && (StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[31 : 2] == StoreBufferPlugin_logic_slots_0_addr[31 : 2]));
  assign when_StoreBufferPlugin_l640_12 = ((StoreBufferPlugin_logic_slots_0_be[0] && StoreBufferPlugin_logic_forwardingLogic_loadMask[0]) && (! _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[0]));
  assign when_StoreBufferPlugin_l640_13 = ((StoreBufferPlugin_logic_slots_0_be[1] && StoreBufferPlugin_logic_forwardingLogic_loadMask[1]) && (! _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[1]));
  assign when_StoreBufferPlugin_l640_14 = ((StoreBufferPlugin_logic_slots_0_be[2] && StoreBufferPlugin_logic_forwardingLogic_loadMask[2]) && (! _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[2]));
  assign when_StoreBufferPlugin_l640_15 = ((StoreBufferPlugin_logic_slots_0_be[3] && StoreBufferPlugin_logic_forwardingLogic_loadMask[3]) && (! _zz_StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask[3]));
  assign StoreBufferPlugin_logic_forwardingLogic_allRequiredBytesHit = ((StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask & StoreBufferPlugin_logic_forwardingLogic_loadMask) == StoreBufferPlugin_logic_forwardingLogic_loadMask);
  assign StoreBufferPlugin_hw_sqQueryPort_rsp_data = StoreBufferPlugin_logic_forwardingLogic_forwardingResult_data;
  assign StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreHasUnknownAddress = 1'b0;
  always @(*) begin
    StoreBufferPlugin_logic_forwardingLogic_dataNotReadyStall = 1'b0;
    if(when_StoreBufferPlugin_l672) begin
      if(when_StoreBufferPlugin_l678) begin
        if(when_StoreBufferPlugin_l681) begin
          StoreBufferPlugin_logic_forwardingLogic_dataNotReadyStall = 1'b1;
        end
      end
    end
    if(when_StoreBufferPlugin_l672_1) begin
      if(when_StoreBufferPlugin_l678_1) begin
        if(when_StoreBufferPlugin_l681_1) begin
          StoreBufferPlugin_logic_forwardingLogic_dataNotReadyStall = 1'b1;
        end
      end
    end
    if(when_StoreBufferPlugin_l672_2) begin
      if(when_StoreBufferPlugin_l678_2) begin
        if(when_StoreBufferPlugin_l681_2) begin
          StoreBufferPlugin_logic_forwardingLogic_dataNotReadyStall = 1'b1;
        end
      end
    end
    if(when_StoreBufferPlugin_l672_3) begin
      if(when_StoreBufferPlugin_l678_3) begin
        if(when_StoreBufferPlugin_l681_3) begin
          StoreBufferPlugin_logic_forwardingLogic_dataNotReadyStall = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_forwardingLogic_hasOlderOverlappingStore = 1'b0;
    if(when_StoreBufferPlugin_l672) begin
      if(when_StoreBufferPlugin_l678) begin
        StoreBufferPlugin_logic_forwardingLogic_hasOlderOverlappingStore = 1'b1;
      end
    end
    if(when_StoreBufferPlugin_l672_1) begin
      if(when_StoreBufferPlugin_l678_1) begin
        StoreBufferPlugin_logic_forwardingLogic_hasOlderOverlappingStore = 1'b1;
      end
    end
    if(when_StoreBufferPlugin_l672_2) begin
      if(when_StoreBufferPlugin_l678_2) begin
        StoreBufferPlugin_logic_forwardingLogic_hasOlderOverlappingStore = 1'b1;
      end
    end
    if(when_StoreBufferPlugin_l672_3) begin
      if(when_StoreBufferPlugin_l678_3) begin
        StoreBufferPlugin_logic_forwardingLogic_hasOlderOverlappingStore = 1'b1;
      end
    end
  end

  assign when_StoreBufferPlugin_l672 = ((StoreBufferPlugin_logic_slots_0_valid && (! StoreBufferPlugin_logic_slots_0_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_0_isFlush));
  assign _zz_when_StoreBufferPlugin_l678 = StoreBufferPlugin_logic_slots_0_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l678_1 = StoreBufferPlugin_logic_slots_0_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l678_2 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l678_3 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l678_4 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[31 : 2];
  assign _zz_when_StoreBufferPlugin_l678_5 = StoreBufferPlugin_logic_slots_0_addr[31 : 2];
  assign when_StoreBufferPlugin_l678 = ((! (((_zz_when_StoreBufferPlugin_l678 == _zz_when_StoreBufferPlugin_l678_2) && (_zz_when_StoreBufferPlugin_l678_3 <= _zz_when_StoreBufferPlugin_l678_1)) || ((_zz_when_StoreBufferPlugin_l678 != _zz_when_StoreBufferPlugin_l678_2) && (_zz_when_StoreBufferPlugin_l678_1 < _zz_when_StoreBufferPlugin_l678_3)))) && (_zz_when_StoreBufferPlugin_l678_4 == _zz_when_StoreBufferPlugin_l678_5));
  assign when_StoreBufferPlugin_l681 = ((StoreBufferPlugin_logic_slots_0_waitRsp || StoreBufferPlugin_logic_slots_0_isWaitingForRefill) || StoreBufferPlugin_logic_slots_0_isWaitingForWb);
  assign when_StoreBufferPlugin_l672_1 = ((StoreBufferPlugin_logic_slots_1_valid && (! StoreBufferPlugin_logic_slots_1_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_1_isFlush));
  assign _zz_when_StoreBufferPlugin_l678_6 = StoreBufferPlugin_logic_slots_1_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l678_7 = StoreBufferPlugin_logic_slots_1_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l678_8 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l678_9 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l678_10 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[31 : 2];
  assign _zz_when_StoreBufferPlugin_l678_11 = StoreBufferPlugin_logic_slots_1_addr[31 : 2];
  assign when_StoreBufferPlugin_l678_1 = ((! (((_zz_when_StoreBufferPlugin_l678_6 == _zz_when_StoreBufferPlugin_l678_8) && (_zz_when_StoreBufferPlugin_l678_9 <= _zz_when_StoreBufferPlugin_l678_7)) || ((_zz_when_StoreBufferPlugin_l678_6 != _zz_when_StoreBufferPlugin_l678_8) && (_zz_when_StoreBufferPlugin_l678_7 < _zz_when_StoreBufferPlugin_l678_9)))) && (_zz_when_StoreBufferPlugin_l678_10 == _zz_when_StoreBufferPlugin_l678_11));
  assign when_StoreBufferPlugin_l681_1 = ((StoreBufferPlugin_logic_slots_1_waitRsp || StoreBufferPlugin_logic_slots_1_isWaitingForRefill) || StoreBufferPlugin_logic_slots_1_isWaitingForWb);
  assign when_StoreBufferPlugin_l672_2 = ((StoreBufferPlugin_logic_slots_2_valid && (! StoreBufferPlugin_logic_slots_2_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_2_isFlush));
  assign _zz_when_StoreBufferPlugin_l678_12 = StoreBufferPlugin_logic_slots_2_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l678_13 = StoreBufferPlugin_logic_slots_2_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l678_14 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l678_15 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l678_16 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[31 : 2];
  assign _zz_when_StoreBufferPlugin_l678_17 = StoreBufferPlugin_logic_slots_2_addr[31 : 2];
  assign when_StoreBufferPlugin_l678_2 = ((! (((_zz_when_StoreBufferPlugin_l678_12 == _zz_when_StoreBufferPlugin_l678_14) && (_zz_when_StoreBufferPlugin_l678_15 <= _zz_when_StoreBufferPlugin_l678_13)) || ((_zz_when_StoreBufferPlugin_l678_12 != _zz_when_StoreBufferPlugin_l678_14) && (_zz_when_StoreBufferPlugin_l678_13 < _zz_when_StoreBufferPlugin_l678_15)))) && (_zz_when_StoreBufferPlugin_l678_16 == _zz_when_StoreBufferPlugin_l678_17));
  assign when_StoreBufferPlugin_l681_2 = ((StoreBufferPlugin_logic_slots_2_waitRsp || StoreBufferPlugin_logic_slots_2_isWaitingForRefill) || StoreBufferPlugin_logic_slots_2_isWaitingForWb);
  assign when_StoreBufferPlugin_l672_3 = ((StoreBufferPlugin_logic_slots_3_valid && (! StoreBufferPlugin_logic_slots_3_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_3_isFlush));
  assign _zz_when_StoreBufferPlugin_l678_18 = StoreBufferPlugin_logic_slots_3_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l678_19 = StoreBufferPlugin_logic_slots_3_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l678_20 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[3];
  assign _zz_when_StoreBufferPlugin_l678_21 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr[2 : 0];
  assign _zz_when_StoreBufferPlugin_l678_22 = StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address[31 : 2];
  assign _zz_when_StoreBufferPlugin_l678_23 = StoreBufferPlugin_logic_slots_3_addr[31 : 2];
  assign when_StoreBufferPlugin_l678_3 = ((! (((_zz_when_StoreBufferPlugin_l678_18 == _zz_when_StoreBufferPlugin_l678_20) && (_zz_when_StoreBufferPlugin_l678_21 <= _zz_when_StoreBufferPlugin_l678_19)) || ((_zz_when_StoreBufferPlugin_l678_18 != _zz_when_StoreBufferPlugin_l678_20) && (_zz_when_StoreBufferPlugin_l678_19 < _zz_when_StoreBufferPlugin_l678_21)))) && (_zz_when_StoreBufferPlugin_l678_22 == _zz_when_StoreBufferPlugin_l678_23));
  assign when_StoreBufferPlugin_l681_3 = ((StoreBufferPlugin_logic_slots_3_waitRsp || StoreBufferPlugin_logic_slots_3_isWaitingForRefill) || StoreBufferPlugin_logic_slots_3_isWaitingForWb);
  assign StoreBufferPlugin_logic_forwardingLogic_insufficientCoverageStall = ((StoreBufferPlugin_hw_sqQueryPort_cmd_valid && StoreBufferPlugin_logic_forwardingLogic_hasOlderOverlappingStore) && (! StoreBufferPlugin_logic_forwardingLogic_allRequiredBytesHit));
  assign StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreDataNotReady = (StoreBufferPlugin_logic_forwardingLogic_dataNotReadyStall || StoreBufferPlugin_logic_forwardingLogic_insufficientCoverageStall);
  assign StoreBufferPlugin_hw_sqQueryPort_rsp_hit = (((StoreBufferPlugin_hw_sqQueryPort_cmd_valid && StoreBufferPlugin_logic_forwardingLogic_allRequiredBytesHit) && (! StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreHasUnknownAddress)) && (! StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreDataNotReady));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_loadQueryBe = 4'b0000;
    case(StoreBufferPlugin_hw_bypassQuerySizeIn)
      MemAccessSize_B : begin
        _zz_StoreBufferPlugin_logic_loadQueryBe = _zz__zz_StoreBufferPlugin_logic_loadQueryBe;
      end
      MemAccessSize_H : begin
        _zz_StoreBufferPlugin_logic_loadQueryBe = _zz__zz_StoreBufferPlugin_logic_loadQueryBe_2[3:0];
      end
      MemAccessSize_W : begin
        _zz_StoreBufferPlugin_logic_loadQueryBe = _zz__zz_StoreBufferPlugin_logic_loadQueryBe_5[3:0];
      end
      default : begin
        _zz_StoreBufferPlugin_logic_loadQueryBe = 4'b1111;
      end
    endcase
  end

  assign _zz_StoreBufferPlugin_logic_loadQueryBe_1 = _zz__zz_StoreBufferPlugin_logic_loadQueryBe_1[1 : 0];
  assign StoreBufferPlugin_logic_loadQueryBe = _zz_StoreBufferPlugin_logic_loadQueryBe;
  assign StoreBufferPlugin_logic_bypassInitial_data = 32'h0;
  assign StoreBufferPlugin_logic_bypassInitial_hitMask = 4'b0000;
  always @(*) begin
    _zz_StoreBufferPlugin_logic_finalBypassResult_data = StoreBufferPlugin_logic_bypassInitial_data;
    if(when_StoreBufferPlugin_l735) begin
      if(when_StoreBufferPlugin_l740) begin
        if(when_StoreBufferPlugin_l742) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data[7 : 0] = StoreBufferPlugin_logic_slots_3_data[7 : 0];
        end
        if(when_StoreBufferPlugin_l742_1) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data[15 : 8] = StoreBufferPlugin_logic_slots_3_data[15 : 8];
        end
        if(when_StoreBufferPlugin_l742_2) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data[23 : 16] = StoreBufferPlugin_logic_slots_3_data[23 : 16];
        end
        if(when_StoreBufferPlugin_l742_3) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data[31 : 24] = StoreBufferPlugin_logic_slots_3_data[31 : 24];
        end
      end
    end
  end

  always @(*) begin
    _zz_when_StoreBufferPlugin_l742 = StoreBufferPlugin_logic_bypassInitial_hitMask;
    if(when_StoreBufferPlugin_l735) begin
      if(when_StoreBufferPlugin_l740) begin
        if(when_StoreBufferPlugin_l742) begin
          _zz_when_StoreBufferPlugin_l742[0] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_1) begin
          _zz_when_StoreBufferPlugin_l742[1] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_2) begin
          _zz_when_StoreBufferPlugin_l742[2] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_3) begin
          _zz_when_StoreBufferPlugin_l742[3] = 1'b1;
        end
      end
    end
  end

  assign when_StoreBufferPlugin_l735 = ((StoreBufferPlugin_logic_slots_3_valid && (! StoreBufferPlugin_logic_slots_3_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_3_isFlush));
  assign when_StoreBufferPlugin_l740 = (StoreBufferPlugin_hw_bypassQueryAddrIn[31 : 2] == StoreBufferPlugin_logic_slots_3_addr[31 : 2]);
  assign when_StoreBufferPlugin_l742 = ((StoreBufferPlugin_logic_slots_3_be[0] && StoreBufferPlugin_logic_loadQueryBe[0]) && (! StoreBufferPlugin_logic_bypassInitial_hitMask[0]));
  assign when_StoreBufferPlugin_l742_1 = ((StoreBufferPlugin_logic_slots_3_be[1] && StoreBufferPlugin_logic_loadQueryBe[1]) && (! StoreBufferPlugin_logic_bypassInitial_hitMask[1]));
  assign when_StoreBufferPlugin_l742_2 = ((StoreBufferPlugin_logic_slots_3_be[2] && StoreBufferPlugin_logic_loadQueryBe[2]) && (! StoreBufferPlugin_logic_bypassInitial_hitMask[2]));
  assign when_StoreBufferPlugin_l742_3 = ((StoreBufferPlugin_logic_slots_3_be[3] && StoreBufferPlugin_logic_loadQueryBe[3]) && (! StoreBufferPlugin_logic_bypassInitial_hitMask[3]));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_finalBypassResult_data_1 = _zz_StoreBufferPlugin_logic_finalBypassResult_data;
    if(when_StoreBufferPlugin_l735_1) begin
      if(when_StoreBufferPlugin_l740_1) begin
        if(when_StoreBufferPlugin_l742_4) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data_1[7 : 0] = StoreBufferPlugin_logic_slots_2_data[7 : 0];
        end
        if(when_StoreBufferPlugin_l742_5) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data_1[15 : 8] = StoreBufferPlugin_logic_slots_2_data[15 : 8];
        end
        if(when_StoreBufferPlugin_l742_6) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data_1[23 : 16] = StoreBufferPlugin_logic_slots_2_data[23 : 16];
        end
        if(when_StoreBufferPlugin_l742_7) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data_1[31 : 24] = StoreBufferPlugin_logic_slots_2_data[31 : 24];
        end
      end
    end
  end

  always @(*) begin
    _zz_when_StoreBufferPlugin_l742_1 = _zz_when_StoreBufferPlugin_l742;
    if(when_StoreBufferPlugin_l735_1) begin
      if(when_StoreBufferPlugin_l740_1) begin
        if(when_StoreBufferPlugin_l742_4) begin
          _zz_when_StoreBufferPlugin_l742_1[0] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_5) begin
          _zz_when_StoreBufferPlugin_l742_1[1] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_6) begin
          _zz_when_StoreBufferPlugin_l742_1[2] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_7) begin
          _zz_when_StoreBufferPlugin_l742_1[3] = 1'b1;
        end
      end
    end
  end

  assign when_StoreBufferPlugin_l735_1 = ((StoreBufferPlugin_logic_slots_2_valid && (! StoreBufferPlugin_logic_slots_2_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_2_isFlush));
  assign when_StoreBufferPlugin_l740_1 = (StoreBufferPlugin_hw_bypassQueryAddrIn[31 : 2] == StoreBufferPlugin_logic_slots_2_addr[31 : 2]);
  assign when_StoreBufferPlugin_l742_4 = ((StoreBufferPlugin_logic_slots_2_be[0] && StoreBufferPlugin_logic_loadQueryBe[0]) && (! _zz_when_StoreBufferPlugin_l742[0]));
  assign when_StoreBufferPlugin_l742_5 = ((StoreBufferPlugin_logic_slots_2_be[1] && StoreBufferPlugin_logic_loadQueryBe[1]) && (! _zz_when_StoreBufferPlugin_l742[1]));
  assign when_StoreBufferPlugin_l742_6 = ((StoreBufferPlugin_logic_slots_2_be[2] && StoreBufferPlugin_logic_loadQueryBe[2]) && (! _zz_when_StoreBufferPlugin_l742[2]));
  assign when_StoreBufferPlugin_l742_7 = ((StoreBufferPlugin_logic_slots_2_be[3] && StoreBufferPlugin_logic_loadQueryBe[3]) && (! _zz_when_StoreBufferPlugin_l742[3]));
  always @(*) begin
    _zz_StoreBufferPlugin_logic_finalBypassResult_data_2 = _zz_StoreBufferPlugin_logic_finalBypassResult_data_1;
    if(when_StoreBufferPlugin_l735_2) begin
      if(when_StoreBufferPlugin_l740_2) begin
        if(when_StoreBufferPlugin_l742_8) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data_2[7 : 0] = StoreBufferPlugin_logic_slots_1_data[7 : 0];
        end
        if(when_StoreBufferPlugin_l742_9) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data_2[15 : 8] = StoreBufferPlugin_logic_slots_1_data[15 : 8];
        end
        if(when_StoreBufferPlugin_l742_10) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data_2[23 : 16] = StoreBufferPlugin_logic_slots_1_data[23 : 16];
        end
        if(when_StoreBufferPlugin_l742_11) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_data_2[31 : 24] = StoreBufferPlugin_logic_slots_1_data[31 : 24];
        end
      end
    end
  end

  always @(*) begin
    _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask = _zz_when_StoreBufferPlugin_l742_1;
    if(when_StoreBufferPlugin_l735_2) begin
      if(when_StoreBufferPlugin_l740_2) begin
        if(when_StoreBufferPlugin_l742_8) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask[0] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_9) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask[1] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_10) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask[2] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_11) begin
          _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask[3] = 1'b1;
        end
      end
    end
  end

  assign when_StoreBufferPlugin_l735_2 = ((StoreBufferPlugin_logic_slots_1_valid && (! StoreBufferPlugin_logic_slots_1_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_1_isFlush));
  assign when_StoreBufferPlugin_l740_2 = (StoreBufferPlugin_hw_bypassQueryAddrIn[31 : 2] == StoreBufferPlugin_logic_slots_1_addr[31 : 2]);
  assign when_StoreBufferPlugin_l742_8 = ((StoreBufferPlugin_logic_slots_1_be[0] && StoreBufferPlugin_logic_loadQueryBe[0]) && (! _zz_when_StoreBufferPlugin_l742_1[0]));
  assign when_StoreBufferPlugin_l742_9 = ((StoreBufferPlugin_logic_slots_1_be[1] && StoreBufferPlugin_logic_loadQueryBe[1]) && (! _zz_when_StoreBufferPlugin_l742_1[1]));
  assign when_StoreBufferPlugin_l742_10 = ((StoreBufferPlugin_logic_slots_1_be[2] && StoreBufferPlugin_logic_loadQueryBe[2]) && (! _zz_when_StoreBufferPlugin_l742_1[2]));
  assign when_StoreBufferPlugin_l742_11 = ((StoreBufferPlugin_logic_slots_1_be[3] && StoreBufferPlugin_logic_loadQueryBe[3]) && (! _zz_when_StoreBufferPlugin_l742_1[3]));
  always @(*) begin
    StoreBufferPlugin_logic_finalBypassResult_data = _zz_StoreBufferPlugin_logic_finalBypassResult_data_2;
    if(when_StoreBufferPlugin_l735_3) begin
      if(when_StoreBufferPlugin_l740_3) begin
        if(when_StoreBufferPlugin_l742_12) begin
          StoreBufferPlugin_logic_finalBypassResult_data[7 : 0] = StoreBufferPlugin_logic_slots_0_data[7 : 0];
        end
        if(when_StoreBufferPlugin_l742_13) begin
          StoreBufferPlugin_logic_finalBypassResult_data[15 : 8] = StoreBufferPlugin_logic_slots_0_data[15 : 8];
        end
        if(when_StoreBufferPlugin_l742_14) begin
          StoreBufferPlugin_logic_finalBypassResult_data[23 : 16] = StoreBufferPlugin_logic_slots_0_data[23 : 16];
        end
        if(when_StoreBufferPlugin_l742_15) begin
          StoreBufferPlugin_logic_finalBypassResult_data[31 : 24] = StoreBufferPlugin_logic_slots_0_data[31 : 24];
        end
      end
    end
  end

  always @(*) begin
    StoreBufferPlugin_logic_finalBypassResult_hitMask = _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask;
    if(when_StoreBufferPlugin_l735_3) begin
      if(when_StoreBufferPlugin_l740_3) begin
        if(when_StoreBufferPlugin_l742_12) begin
          StoreBufferPlugin_logic_finalBypassResult_hitMask[0] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_13) begin
          StoreBufferPlugin_logic_finalBypassResult_hitMask[1] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_14) begin
          StoreBufferPlugin_logic_finalBypassResult_hitMask[2] = 1'b1;
        end
        if(when_StoreBufferPlugin_l742_15) begin
          StoreBufferPlugin_logic_finalBypassResult_hitMask[3] = 1'b1;
        end
      end
    end
  end

  assign when_StoreBufferPlugin_l735_3 = ((StoreBufferPlugin_logic_slots_0_valid && (! StoreBufferPlugin_logic_slots_0_hasEarlyException)) && (! StoreBufferPlugin_logic_slots_0_isFlush));
  assign when_StoreBufferPlugin_l740_3 = (StoreBufferPlugin_hw_bypassQueryAddrIn[31 : 2] == StoreBufferPlugin_logic_slots_0_addr[31 : 2]);
  assign when_StoreBufferPlugin_l742_12 = ((StoreBufferPlugin_logic_slots_0_be[0] && StoreBufferPlugin_logic_loadQueryBe[0]) && (! _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask[0]));
  assign when_StoreBufferPlugin_l742_13 = ((StoreBufferPlugin_logic_slots_0_be[1] && StoreBufferPlugin_logic_loadQueryBe[1]) && (! _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask[1]));
  assign when_StoreBufferPlugin_l742_14 = ((StoreBufferPlugin_logic_slots_0_be[2] && StoreBufferPlugin_logic_loadQueryBe[2]) && (! _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask[2]));
  assign when_StoreBufferPlugin_l742_15 = ((StoreBufferPlugin_logic_slots_0_be[3] && StoreBufferPlugin_logic_loadQueryBe[3]) && (! _zz_StoreBufferPlugin_logic_finalBypassResult_hitMask[3]));
  assign StoreBufferPlugin_logic_overallBypassHit = (|StoreBufferPlugin_logic_finalBypassResult_hitMask);
  assign StoreBufferPlugin_hw_bypassDataOutInst_valid = StoreBufferPlugin_logic_overallBypassHit;
  assign StoreBufferPlugin_hw_bypassDataOutInst_payload_data = StoreBufferPlugin_logic_finalBypassResult_data;
  assign StoreBufferPlugin_hw_bypassDataOutInst_payload_hitMask = StoreBufferPlugin_logic_finalBypassResult_hitMask;
  assign StoreBufferPlugin_hw_bypassDataOutInst_payload_hit = (StoreBufferPlugin_logic_overallBypassHit && (StoreBufferPlugin_logic_finalBypassResult_hitMask == StoreBufferPlugin_logic_loadQueryBe));
  assign LinkerPlugin_logic_allWakeupFlows_0_valid = AluIntEU_AluIntEuPlugin_wakeupSourcePort_valid;
  assign LinkerPlugin_logic_allWakeupFlows_0_payload_physRegIdx = AluIntEU_AluIntEuPlugin_wakeupSourcePort_payload_physRegIdx;
  assign LinkerPlugin_logic_allWakeupFlows_1_valid = MulEU_MulEuPlugin_wakeupSourcePort_valid;
  assign LinkerPlugin_logic_allWakeupFlows_1_payload_physRegIdx = MulEU_MulEuPlugin_wakeupSourcePort_payload_physRegIdx;
  assign LinkerPlugin_logic_allWakeupFlows_2_valid = BranchEU_BranchEuPlugin_wakeupSourcePort_valid;
  assign LinkerPlugin_logic_allWakeupFlows_2_payload_physRegIdx = BranchEU_BranchEuPlugin_wakeupSourcePort_payload_physRegIdx;
  assign LinkerPlugin_logic_allWakeupFlows_3_valid = LsuEU_LsuEuPlugin_wakeupSourcePort_valid;
  assign LinkerPlugin_logic_allWakeupFlows_3_payload_physRegIdx = LsuEU_LsuEuPlugin_wakeupSourcePort_payload_physRegIdx;
  assign LinkerPlugin_logic_allWakeupFlows_4_valid = LoadQueuePlugin_hw_wakeupPort_valid;
  assign LinkerPlugin_logic_allWakeupFlows_4_payload_physRegIdx = LoadQueuePlugin_hw_wakeupPort_payload_physRegIdx;
  always @(*) begin
    BusyTablePlugin_early_setup_clearMask = 64'h0;
    if(CommitPlugin_hw_busyTableClearPort_valid) begin
      BusyTablePlugin_early_setup_clearMask[CommitPlugin_hw_busyTableClearPort_payload] = 1'b1;
    end
    if(AluIntEU_AluIntEuPlugin_setup_clearBusyPort_valid) begin
      BusyTablePlugin_early_setup_clearMask[AluIntEU_AluIntEuPlugin_setup_clearBusyPort_payload] = 1'b1;
    end
    if(MulEU_MulEuPlugin_setup_clearBusyPort_valid) begin
      BusyTablePlugin_early_setup_clearMask[MulEU_MulEuPlugin_setup_clearBusyPort_payload] = 1'b1;
    end
    if(BranchEU_BranchEuPlugin_setup_clearBusyPort_valid) begin
      BusyTablePlugin_early_setup_clearMask[BranchEU_BranchEuPlugin_setup_clearBusyPort_payload] = 1'b1;
    end
    if(LsuEU_LsuEuPlugin_setup_clearBusyPort_valid) begin
      BusyTablePlugin_early_setup_clearMask[LsuEU_LsuEuPlugin_setup_clearBusyPort_payload] = 1'b1;
    end
    if(LoadQueuePlugin_hw_busyTableClearPort_valid) begin
      BusyTablePlugin_early_setup_clearMask[LoadQueuePlugin_hw_busyTableClearPort_payload] = 1'b1;
    end
  end

  always @(*) begin
    BusyTablePlugin_early_setup_setMask = 64'h0;
    if(RenamePlugin_setup_btSetBusyPorts_0_valid) begin
      BusyTablePlugin_early_setup_setMask[RenamePlugin_setup_btSetBusyPorts_0_payload] = 1'b1;
    end
  end

  assign BusyTablePlugin_logic_busyTableNext = ((BusyTablePlugin_early_setup_busyTableReg & (~ BusyTablePlugin_early_setup_clearMask)) | BusyTablePlugin_early_setup_setMask);
  assign BusyTablePlugin_combinationalBusyBits = BusyTablePlugin_logic_busyTableNext;
  assign ICachePlugin_invalidate = 1'b0;
  always @(*) begin
    FetchPipelinePlugin_logic_retryIdCounter_willIncrement = 1'b0;
    if(FetchPipelinePlugin_logic_s4_logic_backpressureRedo) begin
      if(when_FetchPipelinePlugin2_l442) begin
        FetchPipelinePlugin_logic_retryIdCounter_willIncrement = 1'b1;
      end
    end
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l458) begin
          FetchPipelinePlugin_logic_retryIdCounter_willIncrement = 1'b1;
        end
      end
    end
  end

  assign FetchPipelinePlugin_logic_retryIdCounter_willClear = 1'b0;
  assign FetchPipelinePlugin_logic_retryIdCounter_willOverflowIfInc = (FetchPipelinePlugin_logic_retryIdCounter_value == 2'b11);
  assign FetchPipelinePlugin_logic_retryIdCounter_willOverflow = (FetchPipelinePlugin_logic_retryIdCounter_willOverflowIfInc && FetchPipelinePlugin_logic_retryIdCounter_willIncrement);
  always @(*) begin
    if(FetchPipelinePlugin_logic_retryIdCounter_willOverflow) begin
      FetchPipelinePlugin_logic_retryIdCounter_valueNext = 2'b01;
    end else begin
      FetchPipelinePlugin_logic_retryIdCounter_valueNext = (FetchPipelinePlugin_logic_retryIdCounter_value + _zz_FetchPipelinePlugin_logic_retryIdCounter_valueNext);
    end
    if(FetchPipelinePlugin_logic_retryIdCounter_willClear) begin
      FetchPipelinePlugin_logic_retryIdCounter_valueNext = 2'b01;
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_doRetryFlush = 1'b0;
    if(FetchPipelinePlugin_logic_s4_logic_backpressureRedo) begin
      if(when_FetchPipelinePlugin2_l442) begin
        FetchPipelinePlugin_logic_doRetryFlush = 1'b1;
      end
    end
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l458) begin
          FetchPipelinePlugin_logic_doRetryFlush = 1'b1;
        end
      end
    end
  end

  assign FetchPipelinePlugin_logic_hardRedirect_valid = (|CommitPlugin_hw_redirectPort_valid);
  assign FetchPipelinePlugin_logic_hardRedirect_payload = CommitPlugin_hw_redirectPort_payload;
  assign FetchPipelinePlugin_doHardRedirect_listening = FetchPipelinePlugin_logic_hardRedirect_valid;
  assign FetchPipelinePlugin_doSoftRedirect_listening = FetchPipelinePlugin_logic_dispatcher_io_softRedirect_valid;
  assign FetchPipelinePlugin_logic_doAnyFlush = (FetchPipelinePlugin_logic_dispatcher_io_softRedirect_valid || FetchPipelinePlugin_logic_hardRedirect_valid);
  assign io_pop_fire = (FetchPipelinePlugin_setup_fetchOutput_io_pop_valid && s0_Decode_ready);
  always @(*) begin
    FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_incrementIt = 1'b0;
    if(ICachePlugin_port_cmd_valid) begin
      FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_decrementIt = 1'b0;
    if(ICachePlugin_port_rsp_valid) begin
      FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_decrementIt = 1'b1;
    end
  end

  assign FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_mayOverflow = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value == 3'b111);
  assign FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_mayUnderflow = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value == 3'b000);
  assign FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willOverflowIfInc = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_mayOverflow && (! FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_decrementIt));
  assign FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willOverflow = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willOverflowIfInc && FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_incrementIt);
  assign FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willUnderflowIfDec = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_mayUnderflow && (! FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_incrementIt));
  assign FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willUnderflow = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_willUnderflowIfDec && FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_decrementIt);
  assign when_Utils_l767 = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_incrementIt && (! FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l767) begin
      FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l769) begin
        FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_finalIncrement = 3'b111;
      end else begin
        FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l769 = ((! FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_incrementIt) && FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_decrementIt);
  assign FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_valueNext = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value + FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_finalIncrement);
  assign when_FetchPipelinePlugin2_l289 = (FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value == 3'b000);
  assign FetchPipelinePlugin_logic_s1_logic_needRedo = (((FetchPipelinePlugin_logic_retryCmd_lock && (FetchPipelinePlugin_logic_retryCmd_id != FetchPipelinePlugin_logic_s1_logic_lastRetryIdReg)) && (! FetchPipelinePlugin_logic_doAnyFlush)) && (! FetchPipelinePlugin_logic_isDrainingCacheRspReg));
  assign FetchPipelinePlugin_logic_s1_logic_rawPcToUse = (FetchPipelinePlugin_logic_s1_logic_needRedo ? FetchPipelinePlugin_logic_retryCmd_pc : FetchPipelinePlugin_logic_s1_logic_fetchPcReg);
  assign s1_PC_Gen_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC = FetchPipelinePlugin_logic_s1_logic_rawPcToUse;
  assign s1_PC_Gen_FetchPipelinePlugin_logic_FetchPipeline_PC = {FetchPipelinePlugin_logic_s1_logic_rawPcToUse[31 : 4],4'b0000};
  assign FetchPipelinePlugin_logic_s1_logic_nextLinePc = (FetchPipelinePlugin_logic_s1_logic_fetchPcReg + 32'h00000010);
  assign _zz_FetchPipelinePlugin_logic_s1_logic_fetchPcReg = ({FetchPipelinePlugin_logic_retryCmd_pc[31 : 4],4'b0000} + 32'h00000010);
  assign s1_PC_Gen_isFiring = (s1_PC_Gen_valid && s1_PC_Gen_ready);
  assign when_FetchPipelinePlugin2_l361 = ((s1_PC_Gen_isFiring && (! FetchPipelinePlugin_logic_retryCmd_lock)) && (! FetchPipelinePlugin_logic_doAnyFlush));
  assign when_FetchPipelinePlugin2_l367 = (s1_PC_Gen_isFiring && FetchPipelinePlugin_logic_s1_logic_needRedo);
  assign FetchPipelinePlugin_logic_s1_logic_fetchDisabled = 1'b0;
  assign s1_PC_Gen_valid = 1'b1;
  assign when_FetchPipelinePlugin2_l380 = ((FetchPipelinePlugin_logic_isDrainingCacheRspReg || FetchPipelinePlugin_logic_s1_logic_fetchDisabled) || (FetchPipelinePlugin_logic_retryCmd_lock && (FetchPipelinePlugin_logic_retryCmd_id == FetchPipelinePlugin_logic_s1_logic_lastRetryIdReg)));
  assign s1_PC_Gen_haltRequest_FetchPipelinePlugin2_l381 = _zz_s1_PC_Gen_haltRequest_FetchPipelinePlugin2_l381;
  assign s2_ICache_Access_isFiring = (s2_ICache_Access_valid && s2_ICache_Access_ready);
  assign ICachePlugin_port_cmd_valid = ((s2_ICache_Access_isFiring && (! FetchPipelinePlugin_logic_isDrainingCacheRspReg)) && (! FetchPipelinePlugin_logic_doAnyFlush));
  assign FetchPipelinePlugin_logic_s2_logic_cmdPayload_address = s2_ICache_Access_FetchPipelinePlugin_logic_FetchPipeline_PC;
  assign FetchPipelinePlugin_logic_s2_logic_cmdPayload_transactionId = _zz_FetchPipelinePlugin_logic_s2_logic_cmdPayload_transactionId[7:0];
  assign ICachePlugin_port_cmd_payload_address = FetchPipelinePlugin_logic_s2_logic_cmdPayload_address;
  assign ICachePlugin_port_cmd_payload_transactionId = FetchPipelinePlugin_logic_s2_logic_cmdPayload_transactionId;
  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_valid = 1'b0;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_pc = s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_0 = ICachePlugin_port_rsp_payload_instructions_0;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_1 = ICachePlugin_port_rsp_payload_instructions_1;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_2 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_2 = ICachePlugin_port_rsp_payload_instructions_2;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_3 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_instructions_3 = ICachePlugin_port_rsp_payload_instructions_3;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isBranch = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isBranch = _zz_io_push_payload_predecodeInfos_0_isBranch;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isJump = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isJump = FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isJump;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isDirectJump = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isDirectJump = FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isDirectJump;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_jumpOffset = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_jumpOffset = FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_jumpOffset;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isIdle = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_0_isIdle = FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isIdle;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isBranch = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isBranch = _zz_io_push_payload_predecodeInfos_1_isBranch;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isJump = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isJump = FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isJump;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isDirectJump = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isDirectJump = FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isDirectJump;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_jumpOffset = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_jumpOffset = FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_jumpOffset;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isIdle = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_1_isIdle = FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isIdle;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isBranch = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isBranch = _zz_io_push_payload_predecodeInfos_2_isBranch;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isJump = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isJump = FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isJump;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isDirectJump = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isDirectJump = FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isDirectJump;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_jumpOffset = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_jumpOffset = FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_jumpOffset;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isIdle = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_2_isIdle = FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isIdle;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isBranch = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isBranch = _zz_io_push_payload_predecodeInfos_3_isBranch;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isJump = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isJump = FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isJump;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isDirectJump = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isDirectJump = FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isDirectJump;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_jumpOffset = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_jumpOffset = FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_jumpOffset;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isIdle = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_predecodeInfos_3_isIdle = FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isIdle;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_branchMask = 4'bxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_branchMask = {_zz_io_push_payload_predecodeInfos_0_isBranch,{_zz_io_push_payload_predecodeInfos_1_isBranch,{_zz_io_push_payload_predecodeInfos_2_isBranch,_zz_io_push_payload_predecodeInfos_3_isBranch}}};
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_fault = 1'bx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_fault = (! ICachePlugin_port_rsp_payload_wasHit);
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_numValidInstructions = 3'bxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_numValidInstructions = _zz_io_push_payload_numValidInstructions;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_startInstructionIndex = 2'bxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_payload_startInstructionIndex = _zz_io_push_payload_startInstructionIndex;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_instruction = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_instruction = ICachePlugin_port_rsp_payload_instructions_0;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_instruction = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_instruction = ICachePlugin_port_rsp_payload_instructions_1;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_instruction = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_instruction = ICachePlugin_port_rsp_payload_instructions_2;
        end
      end
    end
  end

  always @(*) begin
    FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_instruction = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
      if(!ICachePlugin_port_rsp_payload_redo) begin
        if(when_FetchPipelinePlugin2_l481) begin
          FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_instruction = ICachePlugin_port_rsp_payload_instructions_3;
        end
      end
    end
  end

  assign s4_Predecode_isFiring = (s4_Predecode_valid && s4_Predecode_ready);
  assign FetchPipelinePlugin_logic_s4_logic_handleRsp = (((s4_Predecode_isFiring && ICachePlugin_port_rsp_valid) && (! FetchPipelinePlugin_logic_isDrainingCacheRspReg)) && (! FetchPipelinePlugin_logic_doAnyFlush));
  assign FetchPipelinePlugin_logic_s4_logic_hasHigherPriorityStuff = (FetchPipelinePlugin_logic_doAnyFlush || FetchPipelinePlugin_logic_isDrainingCacheRspReg);
  assign FetchPipelinePlugin_logic_s4_logic_backpressureRedo = ((((((! s4_Predecode_isFiring) && ICachePlugin_port_rsp_valid) && ICachePlugin_port_rsp_payload_wasHit) && (! FetchPipelinePlugin_logic_isDrainingCacheRspReg)) && (! FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_ready)) && (! FetchPipelinePlugin_logic_s4_logic_hasHigherPriorityStuff));
  assign when_FetchPipelinePlugin2_l442 = (! FetchPipelinePlugin_logic_retryCmd_lock);
  assign _zz_70 = (s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC >>> 3'd4);
  assign when_FetchPipelinePlugin2_l458 = (((! FetchPipelinePlugin_logic_retryCmd_lock) || (FetchPipelinePlugin_logic_retryCmd_lock && ({s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC[31 : 4],4'b0000} == {FetchPipelinePlugin_logic_retryCmd_pc[31 : 4],4'b0000}))) && (! FetchPipelinePlugin_logic_s4_logic_hasHigherPriorityStuff));
  assign when_FetchPipelinePlugin2_l467 = (FetchPipelinePlugin_logic_retryCmd_lock && ({s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC[31 : 4],4'b0000} != {FetchPipelinePlugin_logic_retryCmd_pc[31 : 4],4'b0000}));
  assign when_FetchPipelinePlugin2_l476 = (FetchPipelinePlugin_logic_retryCmd_lock && ({s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC[31 : 4],4'b0000} == {FetchPipelinePlugin_logic_retryCmd_pc[31 : 4],4'b0000}));
  assign when_FetchPipelinePlugin2_l481 = ((! FetchPipelinePlugin_logic_retryCmd_lock) || ({s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC[31 : 4],4'b0000} == {FetchPipelinePlugin_logic_retryCmd_pc[31 : 4],4'b0000}));
  assign _zz_io_push_payload_numValidInstructions_1 = (s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC - s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC);
  assign _zz_io_push_payload_numValidInstructions_2 = (_zz_io_push_payload_numValidInstructions_1[3 : 0] >>> 2'd2);
  assign _zz_io_push_payload_startInstructionIndex = _zz_io_push_payload_numValidInstructions_2;
  assign _zz_io_push_payload_predecodeInfos_0_isBranch = FetchPipelinePlugin_logic_s4_logic_predecoders_0_io_predecodeInfo_isBranch;
  assign _zz_io_push_payload_predecodeInfos_1_isBranch = FetchPipelinePlugin_logic_s4_logic_predecoders_1_io_predecodeInfo_isBranch;
  assign _zz_io_push_payload_predecodeInfos_2_isBranch = FetchPipelinePlugin_logic_s4_logic_predecoders_2_io_predecodeInfo_isBranch;
  assign _zz_io_push_payload_predecodeInfos_3_isBranch = FetchPipelinePlugin_logic_s4_logic_predecoders_3_io_predecodeInfo_isBranch;
  assign _zz_io_push_payload_numValidInstructions = (3'b100 - _zz__zz_io_push_payload_numValidInstructions);
  assign s4_Predecode_haltRequest_FetchPipelinePlugin2_l505 = (! FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_ready);
  assign io_push_fire = (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_valid && FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_push_ready);
  assign FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_ready = (FetchPipelinePlugin_logic_dispatcher_io_fetchGroupIn_ready && (! FetchPipelinePlugin_logic_doAnyFlush));
  assign BpuPipelinePlugin_queryPortIn_valid = FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_valid;
  assign BpuPipelinePlugin_queryPortIn_payload_pc = FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_payload_pc;
  assign BpuPipelinePlugin_queryPortIn_payload_transactionId = FetchPipelinePlugin_logic_dispatcher_io_bpuQuery_payload_transactionId;
  assign io_fetchGroupIn_fire = (FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_valid && FetchPipelinePlugin_logic_dispatcher_io_fetchGroupIn_ready);
  assign _zz_71 = _zz__zz_71;
  assign _zz_s2_ICache_Access_isFlushingRoot = (FetchPipelinePlugin_logic_hardRedirect_valid || FetchPipelinePlugin_logic_doRetryFlush);
  assign _zz_s3_ICache_Wait_isFlushingRoot = (FetchPipelinePlugin_logic_hardRedirect_valid || FetchPipelinePlugin_logic_doRetryFlush);
  assign FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_flush = (FetchPipelinePlugin_logic_doAnyFlush || FetchPipelinePlugin_logic_isDrainingCacheRspReg);
  assign s3_ICache_Wait_isFlushed = _zz_s3_ICache_Wait_isFlushingRoot;
  assign s4_Predecode_isFlushed = FetchPipelinePlugin_logic_hardRedirect_valid;
  assign when_Connection_l66_12 = (|{FetchPipelinePlugin_logic_hardRedirect_valid,_zz_s2_ICache_Access_isFlushingRoot});
  assign s2_ICache_Access_isFlushed = when_Connection_l66_12;
  assign s1_PC_Gen_isFlushed = (|{when_Connection_l66_12,FetchPipelinePlugin_logic_hardRedirect_valid});
  assign s1_PC_Gen_isFlushingRoot = (|FetchPipelinePlugin_logic_hardRedirect_valid);
  assign s2_ICache_Access_isFlushingRoot = (|_zz_s2_ICache_Access_isFlushingRoot);
  assign s3_ICache_Wait_isFlushingRoot = (|_zz_s3_ICache_Wait_isFlushingRoot);
  assign s4_Predecode_isFlushingRoot = (|FetchPipelinePlugin_logic_hardRedirect_valid);
  always @(*) begin
    _zz_s2_ICache_Access_valid = s1_PC_Gen_valid;
    if(s1_PC_Gen_isFlushingRoot) begin
      _zz_s2_ICache_Access_valid = 1'b0;
    end
    if(when_Pipeline_l282_2) begin
      _zz_s2_ICache_Access_valid = 1'b0;
    end
  end

  always @(*) begin
    s1_PC_Gen_ready = s1_PC_Gen_ready_output;
    if(when_Pipeline_l282_2) begin
      s1_PC_Gen_ready = 1'b0;
    end
  end

  assign when_Pipeline_l282_2 = (|s1_PC_Gen_haltRequest_FetchPipelinePlugin2_l381);
  always @(*) begin
    _zz_s4_Predecode_valid = s2_ICache_Access_valid;
    if(s2_ICache_Access_isFlushingRoot) begin
      _zz_s4_Predecode_valid = 1'b0;
    end
  end

  assign s2_ICache_Access_ready = s2_ICache_Access_ready_output;
  always @(*) begin
    s4_Predecode_ready = 1'b1;
    if(when_Pipeline_l282_3) begin
      s4_Predecode_ready = 1'b0;
    end
  end

  assign when_Pipeline_l282_3 = (|s4_Predecode_haltRequest_FetchPipelinePlugin2_l505);
  always @(*) begin
    s1_PC_Gen_ready_output = s2_ICache_Access_ready;
    if(when_Connection_l74_3) begin
      s1_PC_Gen_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_3 = (! s2_ICache_Access_valid);
  always @(*) begin
    s2_ICache_Access_ready_output = s4_Predecode_ready;
    if(when_Connection_l74_4) begin
      s2_ICache_Access_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_4 = (! s4_Predecode_valid);
  assign DataCachePlugin_logic_load_hits = LoadQueuePlugin_hw_dCacheLoadPort_cmd_valid;
  assign DataCachePlugin_logic_load_hit = (|DataCachePlugin_logic_load_hits);
  assign DataCachePlugin_logic_load_hits_bools_0 = DataCachePlugin_logic_load_hits[0];
  assign _zz_DataCachePlugin_logic_load_oh[0] = (DataCachePlugin_logic_load_hits_bools_0 && (! 1'b0));
  assign DataCachePlugin_logic_load_oh = _zz_DataCachePlugin_logic_load_oh;
  assign _zz_DataCachePlugin_logic_load_ohHistory_0 = DataCachePlugin_logic_load_oh;
  assign DataCachePlugin_logic_load_ohHistory_0 = _zz_DataCachePlugin_logic_load_ohHistory_0;
  assign DataCachePlugin_logic_load_ohHistory_1 = _zz_DataCachePlugin_logic_load_ohHistory_1;
  assign DataCachePlugin_logic_load_ohHistory_2 = _zz_DataCachePlugin_logic_load_ohHistory_2;
  assign LoadQueuePlugin_hw_dCacheLoadPort_cmd_ready = DataCachePlugin_logic_load_oh[0];
  assign LoadQueuePlugin_hw_dCacheLoadPort_rsp_valid = (DataCachePlugin_setup_cache_io_load_rsp_valid && DataCachePlugin_logic_load_ohHistory_2[0]);
  assign LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_data = DataCachePlugin_setup_cache_io_load_rsp_payload_data;
  assign LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_fault = DataCachePlugin_setup_cache_io_load_rsp_payload_fault;
  assign LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_redo = DataCachePlugin_setup_cache_io_load_rsp_payload_redo;
  assign LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_refillSlot = DataCachePlugin_setup_cache_io_load_rsp_payload_refillSlot;
  assign LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_refillSlotAny = DataCachePlugin_setup_cache_io_load_rsp_payload_refillSlotAny;
  assign LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_id = DataCachePlugin_setup_cache_io_load_rsp_payload_id;
  assign StoreBufferPlugin_hw_dCacheStorePort_cmd_ready = DataCachePlugin_setup_cache_io_store_cmd_ready;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_valid = DataCachePlugin_setup_cache_io_store_rsp_valid;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_fault = DataCachePlugin_setup_cache_io_store_rsp_payload_fault;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_redo = DataCachePlugin_setup_cache_io_store_rsp_payload_redo;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_refillSlot = DataCachePlugin_setup_cache_io_store_rsp_payload_refillSlot;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_refillSlotAny = DataCachePlugin_setup_cache_io_store_rsp_payload_refillSlotAny;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_flush = DataCachePlugin_setup_cache_io_store_rsp_payload_flush;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_prefetch = DataCachePlugin_setup_cache_io_store_rsp_payload_prefetch;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_address = DataCachePlugin_setup_cache_io_store_rsp_payload_address;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_io = DataCachePlugin_setup_cache_io_store_rsp_payload_io;
  assign StoreBufferPlugin_hw_dCacheStorePort_rsp_payload_id = DataCachePlugin_setup_cache_io_store_rsp_payload_id;
  assign ROBPlugin_aggregatedFlushSignal_valid = CommitPlugin_hw_robFlushPort_valid;
  always @(*) begin
    _zz_ROBPlugin_aggregatedFlushSignal_payload_reason = (2'bxx);
    if(CommitPlugin_hw_robFlushPort_valid) begin
      _zz_ROBPlugin_aggregatedFlushSignal_payload_reason = CommitPlugin_hw_robFlushPort_payload_reason;
    end
  end

  always @(*) begin
    _zz_ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr = 4'bxxxx;
    if(CommitPlugin_hw_robFlushPort_valid) begin
      _zz_ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr = CommitPlugin_hw_robFlushPort_payload_targetRobPtr;
    end
  end

  assign ROBPlugin_aggregatedFlushSignal_payload_reason = _zz_ROBPlugin_aggregatedFlushSignal_payload_reason;
  assign ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr = _zz_ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr;
  assign CoreMemSysPlugin_logic_readBridges_0_io_gmbIn_read_rsp_ready = ((LoadQueuePlugin_logic_loadQueue_slots_0_valid && LoadQueuePlugin_logic_loadQueue_slots_0_isIO) && LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp);
  assign CoreMemSysPlugin_logic_roMasters_0_ar_valid = ICachePlugin_axiMaster_ar_valid;
  assign ICachePlugin_axiMaster_ar_ready = CoreMemSysPlugin_logic_roMasters_0_ar_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_ar_payload_addr = ICachePlugin_axiMaster_ar_payload_addr;
  assign CoreMemSysPlugin_logic_roMasters_0_ar_payload_id = ICachePlugin_axiMaster_ar_payload_id;
  assign CoreMemSysPlugin_logic_roMasters_0_ar_payload_len = ICachePlugin_axiMaster_ar_payload_len;
  assign CoreMemSysPlugin_logic_roMasters_0_ar_payload_size = ICachePlugin_axiMaster_ar_payload_size;
  assign CoreMemSysPlugin_logic_roMasters_0_ar_payload_burst = ICachePlugin_axiMaster_ar_payload_burst;
  assign ICachePlugin_axiMaster_r_valid = CoreMemSysPlugin_logic_roMasters_0_r_valid;
  assign CoreMemSysPlugin_logic_roMasters_0_r_ready = ICachePlugin_axiMaster_r_ready;
  assign ICachePlugin_axiMaster_r_payload_data = CoreMemSysPlugin_logic_roMasters_0_r_payload_data;
  assign ICachePlugin_axiMaster_r_payload_last = CoreMemSysPlugin_logic_roMasters_0_r_payload_last;
  assign ICachePlugin_axiMaster_r_payload_id = CoreMemSysPlugin_logic_roMasters_0_r_payload_id;
  assign ICachePlugin_axiMaster_r_payload_resp = CoreMemSysPlugin_logic_roMasters_0_r_payload_resp;
  assign CoreMemSysPlugin_logic_roMasters_0_aw_valid = 1'b0;
  assign CoreMemSysPlugin_logic_roMasters_0_aw_payload_addr = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  assign CoreMemSysPlugin_logic_roMasters_0_aw_payload_id = 4'bxxxx;
  assign CoreMemSysPlugin_logic_roMasters_0_aw_payload_len = 8'bxxxxxxxx;
  assign CoreMemSysPlugin_logic_roMasters_0_aw_payload_size = 3'bxxx;
  assign CoreMemSysPlugin_logic_roMasters_0_aw_payload_burst = 2'bxx;
  assign CoreMemSysPlugin_logic_roMasters_0_w_valid = 1'b0;
  assign CoreMemSysPlugin_logic_roMasters_0_w_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  assign CoreMemSysPlugin_logic_roMasters_0_w_payload_strb = 4'bxxxx;
  assign CoreMemSysPlugin_logic_roMasters_0_w_payload_last = 1'bx;
  assign CoreMemSysPlugin_logic_roMasters_0_b_ready = 1'b0;
  assign when_CheckpointManagerPlugin_l117 = (CheckpointManagerPlugin_restoreCheckpointTrigger && (! CheckpointManagerPlugin_logic_hasValidCheckpoint));
  assign when_CheckpointManagerPlugin_l121 = (CheckpointManagerPlugin_restoreCheckpointTrigger && CheckpointManagerPlugin_logic_hasValidCheckpoint);
  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_valid = 1'b1;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_0 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_0;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_0 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_1 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_1;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_1 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_2 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_2;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_2 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_3 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_3;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_3 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_4 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_4;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_4 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_5 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_5;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_5 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_6 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_6;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_6 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_7 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_7;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_7 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_8 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_8;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_8 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_9 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_9;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_9 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_10 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_10;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_10 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_11 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_11;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_11 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_12 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_12;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_12 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_13 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_13;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_13 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_14 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_14;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_14 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_15 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_15;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_15 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_16 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_16;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_16 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_17 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_17;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_17 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_18 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_18;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_18 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_19 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_19;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_19 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_20 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_20;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_20 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_21 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_21;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_21 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_22 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_22;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_22 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_23 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_23;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_23 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_24 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_24;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_24 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_25 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_25;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_25 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_26 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_26;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_26 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_27 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_27;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_27 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_28 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_28;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_28 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_29 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_29;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_29 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_30 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_30;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_30 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_31 = CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_31;
    end else begin
      RenameMapTablePlugin_early_setup_rat_io_checkpointRestore_payload_mapping_31 = 6'bxxxxxx;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      SimpleFreeListPlugin_early_setup_freeList_io_recover = 1'b1;
    end else begin
      SimpleFreeListPlugin_early_setup_freeList_io_recover = 1'b0;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      CheckpointManagerPlugin_setup_btRestorePort_valid = 1'b1;
    end else begin
      CheckpointManagerPlugin_setup_btRestorePort_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_CheckpointManagerPlugin_l121) begin
      CheckpointManagerPlugin_setup_btRestorePort_payload_busyBits = CheckpointManagerPlugin_logic_storedBtCheckpoint_busyBits;
    end else begin
      CheckpointManagerPlugin_setup_btRestorePort_payload_busyBits = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    ICachePlugin_logic_tag_write_logic_fsmIsCommitting = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
        ICachePlugin_logic_tag_write_logic_fsmIsCommitting = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_logic_tag_write_logic_f2IsUpdatingLru = 1'b0;
    if(ICachePlugin_logic_pipeline_f2_f2_can_update_lru) begin
      ICachePlugin_logic_tag_write_logic_f2IsUpdatingLru = 1'b1;
    end
  end

  always @(*) begin
    ICachePlugin_logic_tag_write_logic_writeAddress = 7'bxxxxxxx;
    if(ICachePlugin_logic_pipeline_f2_f2_can_update_lru) begin
      ICachePlugin_logic_tag_write_logic_writeAddress = ICachePlugin_logic_pipeline_f2_f2_index;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
        ICachePlugin_logic_tag_write_logic_writeAddress = _zz_ICachePlugin_logic_tag_write_logic_writeAddress;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag = 21'bxxxxxxxxxxxxxxxxxxxxx;
    if(ICachePlugin_logic_pipeline_f2_f2_can_update_lru) begin
      ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag = ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_0_tag;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
        ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag = _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag = 21'bxxxxxxxxxxxxxxxxxxxxx;
    if(ICachePlugin_logic_pipeline_f2_f2_can_update_lru) begin
      ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag = ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_1_tag;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
        ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag = _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_logic_tag_write_logic_writeData_lru = 1'bx;
    if(ICachePlugin_logic_pipeline_f2_f2_can_update_lru) begin
      ICachePlugin_logic_tag_write_logic_writeData_lru = (! ICachePlugin_logic_pipeline_f2_hitWayIdx[0]);
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
        ICachePlugin_logic_tag_write_logic_writeData_lru = (! ICachePlugin_logic_refill_victimWayReg[0]);
      end
      default : begin
      end
    endcase
  end

  assign ICachePlugin_logic_tag_write_logic_writeEnable = (ICachePlugin_logic_tag_write_logic_fsmIsCommitting || ICachePlugin_logic_tag_write_logic_f2IsUpdatingLru);
  assign ICache_F1_Access_valid = ICachePlugin_port_cmd_valid;
  assign ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_address = ICachePlugin_port_cmd_payload_address;
  assign ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_transactionId = ICachePlugin_port_cmd_payload_transactionId;
  assign ICachePlugin_logic_pipeline_f1_f1_index = ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_address[10 : 4];
  assign ICache_F1_Access_isFiring = (ICache_F1_Access_valid && ICache_F1_Access_ready);
  assign ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 = _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0;
  assign ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 = _zz_ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1;
  assign _zz_ICachePlugin_logic_pipeline_f1_metaReadData_lru = ICachePlugin_logic_storage_tagLruRam_spinal_port1;
  assign _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag = _zz_ICachePlugin_logic_pipeline_f1_metaReadData_lru[41 : 0];
  assign ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag = _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag_1[20 : 0];
  assign ICachePlugin_logic_pipeline_f1_metaReadData_ways_1_tag = _zz_ICachePlugin_logic_pipeline_f1_metaReadData_ways_1_tag[20 : 0];
  assign ICachePlugin_logic_pipeline_f1_metaReadData_lru = _zz_ICachePlugin_logic_pipeline_f1_metaReadData_lru[42];
  assign _zz_ICachePlugin_logic_pipeline_f1_dataReadData_0_0 = ICachePlugin_logic_storage_dataRams_0_spinal_port0;
  assign ICachePlugin_logic_pipeline_f1_dataReadData_0_0 = _zz_ICachePlugin_logic_pipeline_f1_dataReadData_0_0[31 : 0];
  assign ICachePlugin_logic_pipeline_f1_dataReadData_0_1 = _zz_ICachePlugin_logic_pipeline_f1_dataReadData_0_0[63 : 32];
  assign ICachePlugin_logic_pipeline_f1_dataReadData_0_2 = _zz_ICachePlugin_logic_pipeline_f1_dataReadData_0_0[95 : 64];
  assign ICachePlugin_logic_pipeline_f1_dataReadData_0_3 = _zz_ICachePlugin_logic_pipeline_f1_dataReadData_0_0[127 : 96];
  assign _zz_ICachePlugin_logic_pipeline_f1_dataReadData_1_0 = ICachePlugin_logic_storage_dataRams_1_spinal_port0;
  assign ICachePlugin_logic_pipeline_f1_dataReadData_1_0 = _zz_ICachePlugin_logic_pipeline_f1_dataReadData_1_0[31 : 0];
  assign ICachePlugin_logic_pipeline_f1_dataReadData_1_1 = _zz_ICachePlugin_logic_pipeline_f1_dataReadData_1_0[63 : 32];
  assign ICachePlugin_logic_pipeline_f1_dataReadData_1_2 = _zz_ICachePlugin_logic_pipeline_f1_dataReadData_1_0[95 : 64];
  assign ICachePlugin_logic_pipeline_f1_dataReadData_1_3 = _zz_ICachePlugin_logic_pipeline_f1_dataReadData_1_0[127 : 96];
  assign ICachePlugin_logic_pipeline_f1_writeReadHazard = (ICachePlugin_logic_tag_write_logic_writeEnable && (ICachePlugin_logic_tag_write_logic_writeAddress == ICachePlugin_logic_pipeline_f1_f1_index));
  assign ICache_F1_Access_ICachePlugin_logic_pipeline_F2_USE_FORWARDED_META = ICachePlugin_logic_pipeline_f1_writeReadHazard;
  assign ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_0_tag = ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag;
  assign ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_1_tag = ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag;
  assign ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_lru = ICachePlugin_logic_tag_write_logic_writeData_lru;
  assign ICachePlugin_logic_pipeline_f2_f2_index = ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_address[10 : 4];
  assign ICachePlugin_logic_pipeline_f2_f2_tag = ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_address[31 : 11];
  assign ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_0_tag = (ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_USE_FORWARDED_META ? ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_0_tag : ICachePlugin_logic_pipeline_f1_metaReadData_ways_0_tag);
  assign ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_1_tag = (ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_USE_FORWARDED_META ? ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_1_tag : ICachePlugin_logic_pipeline_f1_metaReadData_ways_1_tag);
  assign ICachePlugin_logic_pipeline_f2_f2_metaLine_lru = (ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_USE_FORWARDED_META ? ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_lru : ICachePlugin_logic_pipeline_f1_metaReadData_lru);
  assign ICachePlugin_logic_pipeline_f2_hit_ways_0 = (ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 && (ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_0_tag == ICachePlugin_logic_pipeline_f2_f2_tag));
  assign ICachePlugin_logic_pipeline_f2_hit_ways_1 = (ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 && (ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_1_tag == ICachePlugin_logic_pipeline_f2_f2_tag));
  assign ICachePlugin_logic_pipeline_f2_isHit = (|{ICachePlugin_logic_pipeline_f2_hit_ways_1,ICachePlugin_logic_pipeline_f2_hit_ways_0});
  assign ICachePlugin_logic_pipeline_f2_hitWayData_0 = (ICachePlugin_logic_pipeline_f2_hit_ways_0 ? ICachePlugin_logic_pipeline_f1_dataReadData_0_0 : ICachePlugin_logic_pipeline_f1_dataReadData_1_0);
  assign ICachePlugin_logic_pipeline_f2_hitWayData_1 = (ICachePlugin_logic_pipeline_f2_hit_ways_0 ? ICachePlugin_logic_pipeline_f1_dataReadData_0_1 : ICachePlugin_logic_pipeline_f1_dataReadData_1_1);
  assign ICachePlugin_logic_pipeline_f2_hitWayData_2 = (ICachePlugin_logic_pipeline_f2_hit_ways_0 ? ICachePlugin_logic_pipeline_f1_dataReadData_0_2 : ICachePlugin_logic_pipeline_f1_dataReadData_1_2);
  assign ICachePlugin_logic_pipeline_f2_hitWayData_3 = (ICachePlugin_logic_pipeline_f2_hit_ways_0 ? ICachePlugin_logic_pipeline_f1_dataReadData_0_3 : ICachePlugin_logic_pipeline_f1_dataReadData_1_3);
  assign _zz_ICachePlugin_logic_pipeline_f2_hitWayIdx = _zz__zz_ICachePlugin_logic_pipeline_f2_hitWayIdx[1];
  assign ICachePlugin_logic_pipeline_f2_hitWayIdx = _zz_ICachePlugin_logic_pipeline_f2_hitWayIdx;
  assign ICache_F2_HitCheck_isFiring = (ICache_F2_HitCheck_valid && ICache_F2_HitCheck_ready);
  assign ICachePlugin_logic_pipeline_f2_f2_can_update_lru = (ICache_F2_HitCheck_isFiring && ICachePlugin_logic_pipeline_f2_isHit);
  always @(*) begin
    ICachePlugin_port_rsp_valid = 1'b0;
    if(ICache_F2_HitCheck_valid) begin
      ICachePlugin_port_rsp_valid = 1'b1;
    end
  end

  always @(*) begin
    ICachePlugin_port_rsp_payload_transactionId = 8'bxxxxxxxx;
    if(ICache_F2_HitCheck_valid) begin
      ICachePlugin_port_rsp_payload_transactionId = ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_transactionId;
    end
  end

  always @(*) begin
    ICachePlugin_port_rsp_payload_instructions_0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(ICache_F2_HitCheck_valid) begin
      if(ICachePlugin_logic_pipeline_f2_isHit) begin
        ICachePlugin_port_rsp_payload_instructions_0 = ICachePlugin_logic_pipeline_f2_hitWayData_0;
      end else begin
        ICachePlugin_port_rsp_payload_instructions_0 = 32'h0;
      end
    end
  end

  always @(*) begin
    ICachePlugin_port_rsp_payload_instructions_1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(ICache_F2_HitCheck_valid) begin
      if(ICachePlugin_logic_pipeline_f2_isHit) begin
        ICachePlugin_port_rsp_payload_instructions_1 = ICachePlugin_logic_pipeline_f2_hitWayData_1;
      end else begin
        ICachePlugin_port_rsp_payload_instructions_1 = 32'h0;
      end
    end
  end

  always @(*) begin
    ICachePlugin_port_rsp_payload_instructions_2 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(ICache_F2_HitCheck_valid) begin
      if(ICachePlugin_logic_pipeline_f2_isHit) begin
        ICachePlugin_port_rsp_payload_instructions_2 = ICachePlugin_logic_pipeline_f2_hitWayData_2;
      end else begin
        ICachePlugin_port_rsp_payload_instructions_2 = 32'h0;
      end
    end
  end

  always @(*) begin
    ICachePlugin_port_rsp_payload_instructions_3 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(ICache_F2_HitCheck_valid) begin
      if(ICachePlugin_logic_pipeline_f2_isHit) begin
        ICachePlugin_port_rsp_payload_instructions_3 = ICachePlugin_logic_pipeline_f2_hitWayData_3;
      end else begin
        ICachePlugin_port_rsp_payload_instructions_3 = 32'h0;
      end
    end
  end

  always @(*) begin
    ICachePlugin_port_rsp_payload_wasHit = 1'bx;
    if(ICache_F2_HitCheck_valid) begin
      ICachePlugin_port_rsp_payload_wasHit = ICachePlugin_logic_pipeline_f2_isHit;
    end
  end

  always @(*) begin
    ICachePlugin_port_rsp_payload_redo = 1'bx;
    if(ICache_F2_HitCheck_valid) begin
      if(ICachePlugin_logic_pipeline_f2_isHit) begin
        ICachePlugin_port_rsp_payload_redo = 1'b0;
      end else begin
        ICachePlugin_port_rsp_payload_redo = 1'b1;
      end
    end
  end

  always @(*) begin
    ICachePlugin_axiMaster_ar_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
        ICachePlugin_axiMaster_ar_valid = 1'b1;
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_axiMaster_ar_payload_addr = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
        ICachePlugin_axiMaster_ar_payload_addr = ICachePlugin_logic_refill_refillCmdReg_address;
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign ICachePlugin_axiMaster_ar_payload_id = 4'bxxxx;
  always @(*) begin
    ICachePlugin_axiMaster_ar_payload_len = 8'bxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
        ICachePlugin_axiMaster_ar_payload_len = 8'h03;
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_axiMaster_ar_payload_size = 3'bxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
        ICachePlugin_axiMaster_ar_payload_size = 3'b010;
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_axiMaster_ar_payload_burst = 2'bxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
        ICachePlugin_axiMaster_ar_payload_burst = 2'b01;
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_axiMaster_r_ready = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
        ICachePlugin_axiMaster_r_ready = 1'b1;
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_logic_refill_refillCounter_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
        if(ICachePlugin_axiMaster_r_fire) begin
          ICachePlugin_logic_refill_refillCounter_willIncrement = 1'b1;
        end
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ICachePlugin_logic_refill_refillCounter_willClear = 1'b0;
    if(ICachePlugin_logic_refill_fsm_onEntry_SEND_REQ) begin
      ICachePlugin_logic_refill_refillCounter_willClear = 1'b1;
    end
  end

  assign ICachePlugin_logic_refill_refillCounter_willOverflowIfInc = (ICachePlugin_logic_refill_refillCounter_value == 2'b11);
  assign ICachePlugin_logic_refill_refillCounter_willOverflow = (ICachePlugin_logic_refill_refillCounter_willOverflowIfInc && ICachePlugin_logic_refill_refillCounter_willIncrement);
  always @(*) begin
    ICachePlugin_logic_refill_refillCounter_valueNext = (ICachePlugin_logic_refill_refillCounter_value + _zz_ICachePlugin_logic_refill_refillCounter_valueNext);
    if(ICachePlugin_logic_refill_refillCounter_willClear) begin
      ICachePlugin_logic_refill_refillCounter_valueNext = 2'b00;
    end
  end

  assign ICachePlugin_logic_refill_fsm_wantExit = 1'b0;
  always @(*) begin
    ICachePlugin_logic_refill_fsm_wantStart = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
        ICachePlugin_logic_refill_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign ICachePlugin_logic_refill_fsm_wantKill = 1'b0;
  always @(*) begin
    ICachePlugin_logic_refill_fsm_stateNext = ICachePlugin_logic_refill_fsm_stateReg;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
        if(when_ICachePlugin_l212) begin
          ICachePlugin_logic_refill_fsm_stateNext = ICachePlugin_logic_refill_fsm_SEND_REQ;
        end
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
        if(ICachePlugin_axiMaster_ar_fire) begin
          ICachePlugin_logic_refill_fsm_stateNext = ICachePlugin_logic_refill_fsm_RECEIVE_DATA;
        end
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
        if(ICachePlugin_axiMaster_r_fire) begin
          if(ICachePlugin_axiMaster_r_payload_last) begin
            ICachePlugin_logic_refill_fsm_stateNext = ICachePlugin_logic_refill_fsm_COMMIT;
          end
        end
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
        ICachePlugin_logic_refill_fsm_stateNext = ICachePlugin_logic_refill_fsm_IDLE;
      end
      default : begin
      end
    endcase
    if(ICachePlugin_logic_refill_fsm_wantStart) begin
      ICachePlugin_logic_refill_fsm_stateNext = ICachePlugin_logic_refill_fsm_IDLE;
    end
    if(ICachePlugin_logic_refill_fsm_wantKill) begin
      ICachePlugin_logic_refill_fsm_stateNext = ICachePlugin_logic_refill_fsm_BOOT;
    end
  end

  assign when_ICachePlugin_l212 = (ICache_F2_HitCheck_valid && (! ICachePlugin_logic_pipeline_f2_isHit));
  assign ICachePlugin_axiMaster_ar_fire = (ICachePlugin_axiMaster_ar_valid && ICachePlugin_axiMaster_ar_ready);
  assign ICachePlugin_axiMaster_r_fire = (ICachePlugin_axiMaster_r_valid && ICachePlugin_axiMaster_r_ready);
  assign _zz_78 = ({3'd0,1'b1} <<< ICachePlugin_logic_refill_refillCounter_value);
  assign _zz_ICachePlugin_logic_tag_write_logic_writeAddress = ICachePlugin_logic_refill_refillCmdReg_address[10 : 4];
  assign when_ICachePlugin_l260 = (ICachePlugin_logic_refill_victimWayReg == 1'b0);
  assign when_ICachePlugin_l260_1 = (ICachePlugin_logic_refill_victimWayReg == 1'b1);
  always @(*) begin
    _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag = ICachePlugin_logic_refill_latchedMetaOnMiss_ways_0_tag;
    if(_zz_79[0]) begin
      _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag = _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag_1;
    end
  end

  always @(*) begin
    _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag = ICachePlugin_logic_refill_latchedMetaOnMiss_ways_1_tag;
    if(_zz_79[1]) begin
      _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_1_tag = _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag_1;
    end
  end

  assign _zz_79 = ({1'd0,1'b1} <<< ICachePlugin_logic_refill_victimWayReg);
  assign _zz_ICachePlugin_logic_tag_write_logic_writeData_ways_0_tag_1 = ICachePlugin_logic_refill_refillCmdReg_address[31 : 11];
  assign _zz_80 = ({127'd0,1'b1} <<< _zz_ICachePlugin_logic_tag_write_logic_writeAddress);
  assign _zz_81 = _zz_80[0];
  assign _zz_82 = _zz_80[1];
  assign _zz_83 = _zz_80[2];
  assign _zz_84 = _zz_80[3];
  assign _zz_85 = _zz_80[4];
  assign _zz_86 = _zz_80[5];
  assign _zz_87 = _zz_80[6];
  assign _zz_88 = _zz_80[7];
  assign _zz_89 = _zz_80[8];
  assign _zz_90 = _zz_80[9];
  assign _zz_91 = _zz_80[10];
  assign _zz_92 = _zz_80[11];
  assign _zz_93 = _zz_80[12];
  assign _zz_94 = _zz_80[13];
  assign _zz_95 = _zz_80[14];
  assign _zz_96 = _zz_80[15];
  assign _zz_97 = _zz_80[16];
  assign _zz_98 = _zz_80[17];
  assign _zz_99 = _zz_80[18];
  assign _zz_100 = _zz_80[19];
  assign _zz_101 = _zz_80[20];
  assign _zz_102 = _zz_80[21];
  assign _zz_103 = _zz_80[22];
  assign _zz_104 = _zz_80[23];
  assign _zz_105 = _zz_80[24];
  assign _zz_106 = _zz_80[25];
  assign _zz_107 = _zz_80[26];
  assign _zz_108 = _zz_80[27];
  assign _zz_109 = _zz_80[28];
  assign _zz_110 = _zz_80[29];
  assign _zz_111 = _zz_80[30];
  assign _zz_112 = _zz_80[31];
  assign _zz_113 = _zz_80[32];
  assign _zz_114 = _zz_80[33];
  assign _zz_115 = _zz_80[34];
  assign _zz_116 = _zz_80[35];
  assign _zz_117 = _zz_80[36];
  assign _zz_118 = _zz_80[37];
  assign _zz_119 = _zz_80[38];
  assign _zz_120 = _zz_80[39];
  assign _zz_121 = _zz_80[40];
  assign _zz_122 = _zz_80[41];
  assign _zz_123 = _zz_80[42];
  assign _zz_124 = _zz_80[43];
  assign _zz_125 = _zz_80[44];
  assign _zz_126 = _zz_80[45];
  assign _zz_127 = _zz_80[46];
  assign _zz_128 = _zz_80[47];
  assign _zz_129 = _zz_80[48];
  assign _zz_130 = _zz_80[49];
  assign _zz_131 = _zz_80[50];
  assign _zz_132 = _zz_80[51];
  assign _zz_133 = _zz_80[52];
  assign _zz_134 = _zz_80[53];
  assign _zz_135 = _zz_80[54];
  assign _zz_136 = _zz_80[55];
  assign _zz_137 = _zz_80[56];
  assign _zz_138 = _zz_80[57];
  assign _zz_139 = _zz_80[58];
  assign _zz_140 = _zz_80[59];
  assign _zz_141 = _zz_80[60];
  assign _zz_142 = _zz_80[61];
  assign _zz_143 = _zz_80[62];
  assign _zz_144 = _zz_80[63];
  assign _zz_145 = _zz_80[64];
  assign _zz_146 = _zz_80[65];
  assign _zz_147 = _zz_80[66];
  assign _zz_148 = _zz_80[67];
  assign _zz_149 = _zz_80[68];
  assign _zz_150 = _zz_80[69];
  assign _zz_151 = _zz_80[70];
  assign _zz_152 = _zz_80[71];
  assign _zz_153 = _zz_80[72];
  assign _zz_154 = _zz_80[73];
  assign _zz_155 = _zz_80[74];
  assign _zz_156 = _zz_80[75];
  assign _zz_157 = _zz_80[76];
  assign _zz_158 = _zz_80[77];
  assign _zz_159 = _zz_80[78];
  assign _zz_160 = _zz_80[79];
  assign _zz_161 = _zz_80[80];
  assign _zz_162 = _zz_80[81];
  assign _zz_163 = _zz_80[82];
  assign _zz_164 = _zz_80[83];
  assign _zz_165 = _zz_80[84];
  assign _zz_166 = _zz_80[85];
  assign _zz_167 = _zz_80[86];
  assign _zz_168 = _zz_80[87];
  assign _zz_169 = _zz_80[88];
  assign _zz_170 = _zz_80[89];
  assign _zz_171 = _zz_80[90];
  assign _zz_172 = _zz_80[91];
  assign _zz_173 = _zz_80[92];
  assign _zz_174 = _zz_80[93];
  assign _zz_175 = _zz_80[94];
  assign _zz_176 = _zz_80[95];
  assign _zz_177 = _zz_80[96];
  assign _zz_178 = _zz_80[97];
  assign _zz_179 = _zz_80[98];
  assign _zz_180 = _zz_80[99];
  assign _zz_181 = _zz_80[100];
  assign _zz_182 = _zz_80[101];
  assign _zz_183 = _zz_80[102];
  assign _zz_184 = _zz_80[103];
  assign _zz_185 = _zz_80[104];
  assign _zz_186 = _zz_80[105];
  assign _zz_187 = _zz_80[106];
  assign _zz_188 = _zz_80[107];
  assign _zz_189 = _zz_80[108];
  assign _zz_190 = _zz_80[109];
  assign _zz_191 = _zz_80[110];
  assign _zz_192 = _zz_80[111];
  assign _zz_193 = _zz_80[112];
  assign _zz_194 = _zz_80[113];
  assign _zz_195 = _zz_80[114];
  assign _zz_196 = _zz_80[115];
  assign _zz_197 = _zz_80[116];
  assign _zz_198 = _zz_80[117];
  assign _zz_199 = _zz_80[118];
  assign _zz_200 = _zz_80[119];
  assign _zz_201 = _zz_80[120];
  assign _zz_202 = _zz_80[121];
  assign _zz_203 = _zz_80[122];
  assign _zz_204 = _zz_80[123];
  assign _zz_205 = _zz_80[124];
  assign _zz_206 = _zz_80[125];
  assign _zz_207 = _zz_80[126];
  assign _zz_208 = _zz_80[127];
  assign _zz_209 = ({1'd0,1'b1} <<< ICachePlugin_logic_refill_victimWayReg);
  assign ICachePlugin_logic_refill_fsm_onExit_BOOT = ((! ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_BOOT_OH_ID]) && (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_BOOT_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onExit_IDLE = ((! ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) && (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onExit_SEND_REQ = ((! ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) && (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onExit_RECEIVE_DATA = ((! ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) && (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onExit_COMMIT = ((! ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) && (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onEntry_BOOT = ((ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_BOOT_OH_ID]) && (! ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_BOOT_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onEntry_IDLE = ((ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) && (! ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onEntry_SEND_REQ = ((ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) && (! ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onEntry_RECEIVE_DATA = ((ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) && (! ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]));
  assign ICachePlugin_logic_refill_fsm_onEntry_COMMIT = ((ICachePlugin_logic_refill_fsm_stateNext[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) && (! ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]));
  always @(*) begin
    ICachePlugin_logic_management_sim_fsmStateId = 3'b111;
    if(when_ICachePlugin_l299) begin
      ICachePlugin_logic_management_sim_fsmStateId = 3'b000;
    end
    if(when_ICachePlugin_l300) begin
      ICachePlugin_logic_management_sim_fsmStateId = 3'b001;
    end
    if(when_ICachePlugin_l301) begin
      ICachePlugin_logic_management_sim_fsmStateId = 3'b010;
    end
    if(when_ICachePlugin_l302) begin
      ICachePlugin_logic_management_sim_fsmStateId = 3'b011;
    end
  end

  assign when_ICachePlugin_l299 = (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]);
  assign when_ICachePlugin_l300 = (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]);
  assign when_ICachePlugin_l301 = (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]);
  assign when_ICachePlugin_l302 = (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]);
  assign ICache_F1_Access_ready = 1'b1;
  assign ICache_F2_HitCheck_ready = 1'b1;
  assign BpuPipelinePlugin_logic_s1_read_valid = BpuPipelinePlugin_queryPortIn_valid;
  assign BpuPipelinePlugin_logic_s1_read_Q_PC = BpuPipelinePlugin_queryPortIn_payload_pc;
  assign BpuPipelinePlugin_logic_s1_read_TRANSACTION_ID = BpuPipelinePlugin_queryPortIn_payload_transactionId;
  assign BpuPipelinePlugin_logic_s1_read_isFiring = (BpuPipelinePlugin_logic_s1_read_valid && BpuPipelinePlugin_logic_s1_read_ready);
  assign _zz_210 = BpuPipelinePlugin_logic_s1_read_Q_PC[11 : 2];
  assign _zz_211 = BpuPipelinePlugin_logic_s1_read_Q_PC[9 : 2];
  assign _zz_BpuPipelinePlugin_logic_phtReadData_s1 = BpuPipelinePlugin_logic_s1_read_Q_PC[11 : 2];
  assign BpuPipelinePlugin_logic_phtReadData_s1 = BpuPipelinePlugin_logic_pht_spinal_port0;
  assign _zz_BpuPipelinePlugin_logic_btbReadData_s1_valid = BpuPipelinePlugin_logic_s1_read_Q_PC[9 : 2];
  assign _zz_BpuPipelinePlugin_logic_btbReadData_s1_valid_1 = BpuPipelinePlugin_logic_btb_spinal_port0;
  assign BpuPipelinePlugin_logic_btbReadData_s1_valid = _zz_BpuPipelinePlugin_logic_btbReadData_s1_valid_1[0];
  assign BpuPipelinePlugin_logic_btbReadData_s1_tag = _zz_BpuPipelinePlugin_logic_btbReadData_s1_valid_1[22 : 1];
  assign BpuPipelinePlugin_logic_btbReadData_s1_target = _zz_BpuPipelinePlugin_logic_btbReadData_s1_valid_1[54 : 23];
  assign BpuPipelinePlugin_logic_phtPrediction = BpuPipelinePlugin_logic_phtReadData_s1[1];
  assign BpuPipelinePlugin_logic_btbHit = (BpuPipelinePlugin_logic_btbReadData_s1_valid && (BpuPipelinePlugin_logic_btbReadData_s1_tag == BpuPipelinePlugin_logic_s2_predict_Q_PC[31 : 10]));
  assign BpuPipelinePlugin_logic_s2_predict_IS_TAKEN = (BpuPipelinePlugin_logic_btbHit && BpuPipelinePlugin_logic_phtPrediction);
  assign BpuPipelinePlugin_logic_s2_predict_TARGET_PC = BpuPipelinePlugin_logic_btbReadData_s1_target;
  assign BpuPipelinePlugin_logic_s2_predict_isFiring = (BpuPipelinePlugin_logic_s2_predict_valid && BpuPipelinePlugin_logic_s2_predict_ready);
  assign _zz_214 = (BpuPipelinePlugin_logic_btbReadData_s1_tag == BpuPipelinePlugin_logic_s2_predict_Q_PC[31 : 10]);
  assign BpuPipelinePlugin_logic_u1_read_valid = BpuPipelinePlugin_updatePortIn_valid;
  assign BpuPipelinePlugin_updatePortIn_ready = BpuPipelinePlugin_logic_u1_read_ready;
  assign BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_pc = BpuPipelinePlugin_updatePortIn_payload_pc;
  assign BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_isTaken = BpuPipelinePlugin_updatePortIn_payload_isTaken;
  assign BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_target = BpuPipelinePlugin_updatePortIn_payload_target;
  assign BpuPipelinePlugin_logic_u1_read_isFiring = (BpuPipelinePlugin_logic_u1_read_valid && BpuPipelinePlugin_logic_u1_read_ready);
  assign _zz_BpuPipelinePlugin_logic_oldPhtState_u1 = BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_pc[11 : 2];
  assign BpuPipelinePlugin_logic_oldPhtState_u1 = BpuPipelinePlugin_logic_pht_spinal_port1;
  always @(*) begin
    case(BpuPipelinePlugin_logic_oldPhtState_u1)
      2'b00 : begin
        BpuPipelinePlugin_logic_newPhtState = (BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken ? 2'b01 : 2'b00);
      end
      2'b01 : begin
        BpuPipelinePlugin_logic_newPhtState = (BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken ? 2'b10 : 2'b00);
      end
      2'b10 : begin
        BpuPipelinePlugin_logic_newPhtState = (BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken ? 2'b11 : 2'b01);
      end
      default : begin
        BpuPipelinePlugin_logic_newPhtState = (BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken ? 2'b11 : 2'b10);
      end
    endcase
  end

  assign BpuPipelinePlugin_logic_u2_write_isFiring = (BpuPipelinePlugin_logic_u2_write_valid && BpuPipelinePlugin_logic_u2_write_ready);
  assign BpuPipelinePlugin_responseFlowOut_valid = BpuPipelinePlugin_logic_s2_predict_valid;
  assign BpuPipelinePlugin_responseFlowOut_payload_isTaken = BpuPipelinePlugin_logic_s2_predict_IS_TAKEN;
  assign BpuPipelinePlugin_responseFlowOut_payload_target = BpuPipelinePlugin_logic_s2_predict_TARGET_PC;
  assign BpuPipelinePlugin_responseFlowOut_payload_transactionId = BpuPipelinePlugin_logic_s2_predict_TRANSACTION_ID;
  assign BpuPipelinePlugin_responseFlowOut_payload_qPc = BpuPipelinePlugin_logic_s2_predict_Q_PC;
  assign BpuPipelinePlugin_logic_s1_read_ready = 1'b1;
  assign BpuPipelinePlugin_logic_s2_predict_ready = 1'b1;
  assign BpuPipelinePlugin_logic_u1_read_ready = 1'b1;
  assign BpuPipelinePlugin_logic_u2_write_ready = 1'b1;
  assign io_isram_addr = CoreMemSysPlugin_hw_baseramCtrl_io_ram_addr;
  assign io_isram_din = CoreMemSysPlugin_hw_baseramCtrl_io_ram_data_write;
  assign io_isram_en = (! CoreMemSysPlugin_hw_baseramCtrl_io_ram_ce_n);
  assign io_isram_re = (! CoreMemSysPlugin_hw_baseramCtrl_io_ram_oe_n);
  assign io_isram_we = (! CoreMemSysPlugin_hw_baseramCtrl_io_ram_we_n);
  assign io_isram_wmask = (~ CoreMemSysPlugin_hw_baseramCtrl_io_ram_be_n);
  assign io_dsram_addr = CoreMemSysPlugin_hw_extramCtrl_io_ram_addr;
  assign io_dsram_din = CoreMemSysPlugin_hw_extramCtrl_io_ram_data_write;
  assign io_dsram_en = (! CoreMemSysPlugin_hw_extramCtrl_io_ram_ce_n);
  assign io_dsram_re = (! CoreMemSysPlugin_hw_extramCtrl_io_ram_oe_n);
  assign io_dsram_we = (! CoreMemSysPlugin_hw_extramCtrl_io_ram_we_n);
  assign io_dsram_wmask = (~ CoreMemSysPlugin_hw_extramCtrl_io_ram_be_n);
  assign io_uart_ar_bits_id = {1'd0, _zz_io_uart_ar_bits_id};
  assign io_uart_ar_bits_addr = uartAxi_ar_payload_addr;
  assign io_uart_ar_bits_len = uartAxi_ar_payload_len;
  assign io_uart_ar_bits_size = uartAxi_ar_payload_size;
  assign io_uart_ar_bits_burst = uartAxi_ar_payload_burst;
  assign io_uart_ar_valid = uartAxi_ar_valid;
  assign uartAxi_ar_ready = io_uart_ar_ready;
  assign uartAxi_r_payload_id = _zz_uartAxi_r_payload_id[6:0];
  assign uartAxi_r_payload_resp = io_uart_r_bits_resp;
  assign uartAxi_r_payload_data = io_uart_r_bits_data;
  assign uartAxi_r_payload_last = io_uart_r_bits_last;
  assign uartAxi_r_valid = io_uart_r_valid;
  assign io_uart_r_ready = uartAxi_r_ready;
  assign io_uart_aw_bits_id = {1'd0, _zz_io_uart_aw_bits_id};
  assign io_uart_aw_bits_addr = uartAxi_aw_payload_addr;
  assign io_uart_aw_bits_len = uartAxi_aw_payload_len;
  assign io_uart_aw_bits_size = uartAxi_aw_payload_size;
  assign io_uart_aw_bits_burst = uartAxi_aw_payload_burst;
  assign io_uart_aw_valid = uartAxi_aw_valid;
  assign uartAxi_aw_ready = io_uart_aw_ready;
  assign io_uart_w_bits_data = uartAxi_w_payload_data;
  assign io_uart_w_bits_strb = uartAxi_w_payload_strb;
  assign io_uart_w_bits_last = uartAxi_w_payload_last;
  assign io_uart_w_valid = uartAxi_w_valid;
  assign uartAxi_w_ready = io_uart_w_ready;
  assign uartAxi_b_payload_id = _zz_uartAxi_b_payload_id[6:0];
  assign uartAxi_b_payload_resp = io_uart_b_bits_resp;
  assign uartAxi_b_valid = io_uart_b_valid;
  assign io_uart_b_ready = uartAxi_b_ready;
  assign uartAxi_ar_valid = axi4ReadOnlyArbiter_5_io_output_ar_valid;
  assign uartAxi_ar_payload_addr = axi4ReadOnlyArbiter_5_io_output_ar_payload_addr;
  assign uartAxi_ar_payload_id = axi4ReadOnlyArbiter_5_io_output_ar_payload_id;
  assign uartAxi_ar_payload_len = axi4ReadOnlyArbiter_5_io_output_ar_payload_len;
  assign uartAxi_ar_payload_size = axi4ReadOnlyArbiter_5_io_output_ar_payload_size;
  assign uartAxi_ar_payload_burst = axi4ReadOnlyArbiter_5_io_output_ar_payload_burst;
  assign uartAxi_r_ready = axi4ReadOnlyArbiter_5_io_output_r_ready;
  assign uartAxi_aw_valid = axi4WriteOnlyArbiter_5_io_output_aw_valid;
  assign uartAxi_aw_payload_addr = axi4WriteOnlyArbiter_5_io_output_aw_payload_addr;
  assign uartAxi_aw_payload_id = axi4WriteOnlyArbiter_5_io_output_aw_payload_id;
  assign uartAxi_aw_payload_len = axi4WriteOnlyArbiter_5_io_output_aw_payload_len;
  assign uartAxi_aw_payload_size = axi4WriteOnlyArbiter_5_io_output_aw_payload_size;
  assign uartAxi_aw_payload_burst = axi4WriteOnlyArbiter_5_io_output_aw_payload_burst;
  assign uartAxi_w_valid = axi4WriteOnlyArbiter_5_io_output_w_valid;
  assign uartAxi_w_payload_data = axi4WriteOnlyArbiter_5_io_output_w_payload_data;
  assign uartAxi_w_payload_strb = axi4WriteOnlyArbiter_5_io_output_w_payload_strb;
  assign uartAxi_w_payload_last = axi4WriteOnlyArbiter_5_io_output_w_payload_last;
  assign uartAxi_b_ready = axi4WriteOnlyArbiter_5_io_output_b_ready;
  assign io_axiOut_readOnly_ar_valid = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_valid;
  assign io_axiOut_readOnly_ar_payload_addr = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_addr;
  assign io_axiOut_readOnly_ar_payload_id = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_id;
  assign io_axiOut_readOnly_ar_payload_len = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_len;
  assign io_axiOut_readOnly_ar_payload_size = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_size;
  assign io_axiOut_readOnly_ar_payload_burst = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_ar_payload_burst;
  assign io_axiOut_readOnly_r_ready = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_r_ready;
  assign io_axiOut_writeOnly_aw_valid = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_valid;
  assign io_axiOut_writeOnly_aw_payload_addr = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_addr;
  assign io_axiOut_writeOnly_aw_payload_id = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_id;
  assign io_axiOut_writeOnly_aw_payload_len = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_len;
  assign io_axiOut_writeOnly_aw_payload_size = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_size;
  assign io_axiOut_writeOnly_aw_payload_burst = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_aw_payload_burst;
  assign io_axiOut_writeOnly_w_valid = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_valid;
  assign io_axiOut_writeOnly_w_payload_data = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_data;
  assign io_axiOut_writeOnly_w_payload_strb = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_strb;
  assign io_axiOut_writeOnly_w_payload_last = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_w_payload_last;
  assign io_axiOut_writeOnly_b_ready = CoreMemSysPlugin_logic_writeBridges_0_io_axiOut_b_ready;
  assign io_axiOut_readOnly_ar_valid_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_valid;
  assign io_axiOut_readOnly_ar_payload_addr_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_addr;
  assign io_axiOut_readOnly_ar_payload_id_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_id;
  assign io_axiOut_readOnly_ar_payload_len_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_len;
  assign io_axiOut_readOnly_ar_payload_size_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_size;
  assign io_axiOut_readOnly_ar_payload_burst_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_ar_payload_burst;
  assign io_axiOut_readOnly_r_ready_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_r_ready;
  assign io_axiOut_writeOnly_aw_valid_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_valid;
  assign io_axiOut_writeOnly_aw_payload_addr_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_addr;
  assign io_axiOut_writeOnly_aw_payload_id_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_id;
  assign io_axiOut_writeOnly_aw_payload_len_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_len;
  assign io_axiOut_writeOnly_aw_payload_size_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_size;
  assign io_axiOut_writeOnly_aw_payload_burst_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_aw_payload_burst;
  assign io_axiOut_writeOnly_w_valid_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_valid;
  assign io_axiOut_writeOnly_w_payload_data_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_data;
  assign io_axiOut_writeOnly_w_payload_strb_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_strb;
  assign io_axiOut_writeOnly_w_payload_last_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_w_payload_last;
  assign io_axiOut_writeOnly_b_ready_1 = CoreMemSysPlugin_logic_readBridges_0_io_axiOut_b_ready;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_ar_valid = DataCachePlugin_setup_dcacheMaster_ar_valid;
  assign DataCachePlugin_setup_dcacheMaster_ar_ready = DataCachePlugin_setup_dcacheMaster_readOnly_ar_ready;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_addr = DataCachePlugin_setup_dcacheMaster_ar_payload_addr;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_id = DataCachePlugin_setup_dcacheMaster_ar_payload_id;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_len = DataCachePlugin_setup_dcacheMaster_ar_payload_len;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_size = DataCachePlugin_setup_dcacheMaster_ar_payload_size;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_burst = DataCachePlugin_setup_dcacheMaster_ar_payload_burst;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_ar_payload_prot = DataCachePlugin_setup_dcacheMaster_ar_payload_prot;
  assign DataCachePlugin_setup_dcacheMaster_r_valid = DataCachePlugin_setup_dcacheMaster_readOnly_r_valid;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_r_ready = DataCachePlugin_setup_dcacheMaster_r_ready;
  assign DataCachePlugin_setup_dcacheMaster_r_payload_data = DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_data;
  assign DataCachePlugin_setup_dcacheMaster_r_payload_last = DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_last;
  assign DataCachePlugin_setup_dcacheMaster_r_payload_id = DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_id;
  assign DataCachePlugin_setup_dcacheMaster_r_payload_resp = DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_resp;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_aw_valid = DataCachePlugin_setup_dcacheMaster_aw_valid;
  assign DataCachePlugin_setup_dcacheMaster_aw_ready = DataCachePlugin_setup_dcacheMaster_writeOnly_aw_ready;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_addr = DataCachePlugin_setup_dcacheMaster_aw_payload_addr;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_id = DataCachePlugin_setup_dcacheMaster_aw_payload_id;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_len = DataCachePlugin_setup_dcacheMaster_aw_payload_len;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_size = DataCachePlugin_setup_dcacheMaster_aw_payload_size;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_burst = DataCachePlugin_setup_dcacheMaster_aw_payload_burst;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_aw_payload_prot = DataCachePlugin_setup_dcacheMaster_aw_payload_prot;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_w_valid = DataCachePlugin_setup_dcacheMaster_w_valid;
  assign DataCachePlugin_setup_dcacheMaster_w_ready = DataCachePlugin_setup_dcacheMaster_writeOnly_w_ready;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_data = DataCachePlugin_setup_dcacheMaster_w_payload_data;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_strb = DataCachePlugin_setup_dcacheMaster_w_payload_strb;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_w_payload_last = DataCachePlugin_setup_dcacheMaster_w_payload_last;
  assign DataCachePlugin_setup_dcacheMaster_b_valid = DataCachePlugin_setup_dcacheMaster_writeOnly_b_valid;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_b_ready = DataCachePlugin_setup_dcacheMaster_b_ready;
  assign DataCachePlugin_setup_dcacheMaster_b_payload_id = DataCachePlugin_setup_dcacheMaster_writeOnly_b_payload_id;
  assign DataCachePlugin_setup_dcacheMaster_b_payload_resp = DataCachePlugin_setup_dcacheMaster_writeOnly_b_payload_resp;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_valid = CoreMemSysPlugin_logic_roMasters_0_ar_valid;
  assign CoreMemSysPlugin_logic_roMasters_0_ar_ready = CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_addr = CoreMemSysPlugin_logic_roMasters_0_ar_payload_addr;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_id = CoreMemSysPlugin_logic_roMasters_0_ar_payload_id;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_len = CoreMemSysPlugin_logic_roMasters_0_ar_payload_len;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_size = CoreMemSysPlugin_logic_roMasters_0_ar_payload_size;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_payload_burst = CoreMemSysPlugin_logic_roMasters_0_ar_payload_burst;
  assign CoreMemSysPlugin_logic_roMasters_0_r_valid = CoreMemSysPlugin_logic_roMasters_0_readOnly_r_valid;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_r_ready = CoreMemSysPlugin_logic_roMasters_0_r_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_r_payload_data = CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_data;
  assign CoreMemSysPlugin_logic_roMasters_0_r_payload_last = CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_last;
  assign CoreMemSysPlugin_logic_roMasters_0_r_payload_id = CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_id;
  assign CoreMemSysPlugin_logic_roMasters_0_r_payload_resp = CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_resp;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_valid = CoreMemSysPlugin_logic_roMasters_0_aw_valid;
  assign CoreMemSysPlugin_logic_roMasters_0_aw_ready = CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_addr = CoreMemSysPlugin_logic_roMasters_0_aw_payload_addr;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_id = CoreMemSysPlugin_logic_roMasters_0_aw_payload_id;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_len = CoreMemSysPlugin_logic_roMasters_0_aw_payload_len;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_size = CoreMemSysPlugin_logic_roMasters_0_aw_payload_size;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_payload_burst = CoreMemSysPlugin_logic_roMasters_0_aw_payload_burst;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_valid = CoreMemSysPlugin_logic_roMasters_0_w_valid;
  assign CoreMemSysPlugin_logic_roMasters_0_w_ready = CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_data = CoreMemSysPlugin_logic_roMasters_0_w_payload_data;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_strb = CoreMemSysPlugin_logic_roMasters_0_w_payload_strb;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_payload_last = CoreMemSysPlugin_logic_roMasters_0_w_payload_last;
  assign CoreMemSysPlugin_logic_roMasters_0_b_valid = CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_valid;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_ready = CoreMemSysPlugin_logic_roMasters_0_b_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_b_payload_id = CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_payload_id;
  assign CoreMemSysPlugin_logic_roMasters_0_b_payload_resp = CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_payload_resp;
  assign io_outputs_0_ar_validPipe_fire = (io_outputs_0_ar_validPipe_valid && io_outputs_0_ar_validPipe_ready);
  assign io_outputs_0_ar_validPipe_valid = io_outputs_0_ar_rValid;
  assign io_outputs_0_ar_validPipe_payload_addr = io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_addr;
  assign io_outputs_0_ar_validPipe_payload_id = io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_id;
  assign io_outputs_0_ar_validPipe_payload_len = io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_len;
  assign io_outputs_0_ar_validPipe_payload_size = io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_size;
  assign io_outputs_0_ar_validPipe_payload_burst = io_axiOut_readOnly_decoder_io_outputs_0_ar_payload_burst;
  assign io_outputs_0_ar_validPipe_ready = axi4ReadOnlyArbiter_3_io_inputs_0_ar_ready;
  assign io_axiOut_readOnly_decoder_io_outputs_0_r_payload_id = axi4ReadOnlyArbiter_3_io_inputs_0_r_payload_id[3:0];
  assign io_outputs_1_ar_validPipe_fire = (io_outputs_1_ar_validPipe_valid && io_outputs_1_ar_validPipe_ready);
  assign io_outputs_1_ar_validPipe_valid = io_outputs_1_ar_rValid;
  assign io_outputs_1_ar_validPipe_payload_addr = io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_addr;
  assign io_outputs_1_ar_validPipe_payload_id = io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_id;
  assign io_outputs_1_ar_validPipe_payload_len = io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_len;
  assign io_outputs_1_ar_validPipe_payload_size = io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_size;
  assign io_outputs_1_ar_validPipe_payload_burst = io_axiOut_readOnly_decoder_io_outputs_1_ar_payload_burst;
  assign io_outputs_1_ar_validPipe_ready = axi4ReadOnlyArbiter_4_io_inputs_0_ar_ready;
  assign io_axiOut_readOnly_decoder_io_outputs_1_r_payload_id = axi4ReadOnlyArbiter_4_io_inputs_0_r_payload_id[3:0];
  assign io_outputs_2_ar_validPipe_fire = (io_outputs_2_ar_validPipe_valid && io_outputs_2_ar_validPipe_ready);
  assign io_outputs_2_ar_validPipe_valid = io_outputs_2_ar_rValid;
  assign io_outputs_2_ar_validPipe_payload_addr = io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_addr;
  assign io_outputs_2_ar_validPipe_payload_id = io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_id;
  assign io_outputs_2_ar_validPipe_payload_len = io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_len;
  assign io_outputs_2_ar_validPipe_payload_size = io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_size;
  assign io_outputs_2_ar_validPipe_payload_burst = io_axiOut_readOnly_decoder_io_outputs_2_ar_payload_burst;
  assign io_outputs_2_ar_validPipe_ready = axi4ReadOnlyArbiter_5_io_inputs_0_ar_ready;
  assign io_axiOut_readOnly_decoder_io_outputs_2_r_payload_id = axi4ReadOnlyArbiter_5_io_inputs_0_r_payload_id[3:0];
  assign io_axiOut_readOnly_ar_ready = io_axiOut_readOnly_decoder_io_input_ar_ready;
  assign io_axiOut_readOnly_r_valid = io_axiOut_readOnly_decoder_io_input_r_valid;
  assign io_axiOut_readOnly_r_payload_data = io_axiOut_readOnly_decoder_io_input_r_payload_data;
  assign io_axiOut_readOnly_r_payload_last = io_axiOut_readOnly_decoder_io_input_r_payload_last;
  assign io_axiOut_readOnly_r_payload_id = io_axiOut_readOnly_decoder_io_input_r_payload_id;
  assign io_axiOut_readOnly_r_payload_resp = io_axiOut_readOnly_decoder_io_input_r_payload_resp;
  assign io_outputs_0_aw_validPipe_fire = (io_outputs_0_aw_validPipe_valid && io_outputs_0_aw_validPipe_ready);
  assign io_outputs_0_aw_validPipe_valid = io_outputs_0_aw_rValid;
  assign io_outputs_0_aw_validPipe_payload_addr = io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  assign io_outputs_0_aw_validPipe_payload_id = io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_id;
  assign io_outputs_0_aw_validPipe_payload_len = io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_len;
  assign io_outputs_0_aw_validPipe_payload_size = io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_size;
  assign io_outputs_0_aw_validPipe_payload_burst = io_axiOut_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  assign io_outputs_0_aw_validPipe_ready = axi4WriteOnlyArbiter_3_io_inputs_0_aw_ready;
  assign io_axiOut_writeOnly_decoder_io_outputs_0_b_payload_id = axi4WriteOnlyArbiter_3_io_inputs_0_b_payload_id[3:0];
  assign io_outputs_1_aw_validPipe_fire = (io_outputs_1_aw_validPipe_valid && io_outputs_1_aw_validPipe_ready);
  assign io_outputs_1_aw_validPipe_valid = io_outputs_1_aw_rValid;
  assign io_outputs_1_aw_validPipe_payload_addr = io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_addr;
  assign io_outputs_1_aw_validPipe_payload_id = io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_id;
  assign io_outputs_1_aw_validPipe_payload_len = io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_len;
  assign io_outputs_1_aw_validPipe_payload_size = io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_size;
  assign io_outputs_1_aw_validPipe_payload_burst = io_axiOut_writeOnly_decoder_io_outputs_1_aw_payload_burst;
  assign io_outputs_1_aw_validPipe_ready = axi4WriteOnlyArbiter_4_io_inputs_0_aw_ready;
  assign io_axiOut_writeOnly_decoder_io_outputs_1_b_payload_id = axi4WriteOnlyArbiter_4_io_inputs_0_b_payload_id[3:0];
  assign io_outputs_2_aw_validPipe_fire = (io_outputs_2_aw_validPipe_valid && io_outputs_2_aw_validPipe_ready);
  assign io_outputs_2_aw_validPipe_valid = io_outputs_2_aw_rValid;
  assign io_outputs_2_aw_validPipe_payload_addr = io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_addr;
  assign io_outputs_2_aw_validPipe_payload_id = io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_id;
  assign io_outputs_2_aw_validPipe_payload_len = io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_len;
  assign io_outputs_2_aw_validPipe_payload_size = io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_size;
  assign io_outputs_2_aw_validPipe_payload_burst = io_axiOut_writeOnly_decoder_io_outputs_2_aw_payload_burst;
  assign io_outputs_2_aw_validPipe_ready = axi4WriteOnlyArbiter_5_io_inputs_0_aw_ready;
  assign io_axiOut_writeOnly_decoder_io_outputs_2_b_payload_id = axi4WriteOnlyArbiter_5_io_inputs_0_b_payload_id[3:0];
  assign io_axiOut_writeOnly_aw_ready = io_axiOut_writeOnly_decoder_io_input_aw_ready;
  assign io_axiOut_writeOnly_w_ready = io_axiOut_writeOnly_decoder_io_input_w_ready;
  assign io_axiOut_writeOnly_b_valid = io_axiOut_writeOnly_decoder_io_input_b_valid;
  assign io_axiOut_writeOnly_b_payload_id = io_axiOut_writeOnly_decoder_io_input_b_payload_id;
  assign io_axiOut_writeOnly_b_payload_resp = io_axiOut_writeOnly_decoder_io_input_b_payload_resp;
  assign io_outputs_0_ar_validPipe_fire_1 = (io_outputs_0_ar_validPipe_valid_1 && io_outputs_0_ar_validPipe_ready_1);
  assign io_outputs_0_ar_validPipe_valid_1 = io_outputs_0_ar_rValid_1;
  assign io_outputs_0_ar_validPipe_payload_addr_1 = io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_addr;
  assign io_outputs_0_ar_validPipe_payload_id_1 = io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_id;
  assign io_outputs_0_ar_validPipe_payload_len_1 = io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_len;
  assign io_outputs_0_ar_validPipe_payload_size_1 = io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_size;
  assign io_outputs_0_ar_validPipe_payload_burst_1 = io_axiOut_readOnly_decoder_1_io_outputs_0_ar_payload_burst;
  assign io_outputs_0_ar_validPipe_ready_1 = axi4ReadOnlyArbiter_3_io_inputs_1_ar_ready;
  assign io_axiOut_readOnly_decoder_1_io_outputs_0_r_payload_id = axi4ReadOnlyArbiter_3_io_inputs_1_r_payload_id[3:0];
  assign io_outputs_1_ar_validPipe_fire_1 = (io_outputs_1_ar_validPipe_valid_1 && io_outputs_1_ar_validPipe_ready_1);
  assign io_outputs_1_ar_validPipe_valid_1 = io_outputs_1_ar_rValid_1;
  assign io_outputs_1_ar_validPipe_payload_addr_1 = io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_addr;
  assign io_outputs_1_ar_validPipe_payload_id_1 = io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_id;
  assign io_outputs_1_ar_validPipe_payload_len_1 = io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_len;
  assign io_outputs_1_ar_validPipe_payload_size_1 = io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_size;
  assign io_outputs_1_ar_validPipe_payload_burst_1 = io_axiOut_readOnly_decoder_1_io_outputs_1_ar_payload_burst;
  assign io_outputs_1_ar_validPipe_ready_1 = axi4ReadOnlyArbiter_4_io_inputs_1_ar_ready;
  assign io_axiOut_readOnly_decoder_1_io_outputs_1_r_payload_id = axi4ReadOnlyArbiter_4_io_inputs_1_r_payload_id[3:0];
  assign io_outputs_2_ar_validPipe_fire_1 = (io_outputs_2_ar_validPipe_valid_1 && io_outputs_2_ar_validPipe_ready_1);
  assign io_outputs_2_ar_validPipe_valid_1 = io_outputs_2_ar_rValid_1;
  assign io_outputs_2_ar_validPipe_payload_addr_1 = io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_addr;
  assign io_outputs_2_ar_validPipe_payload_id_1 = io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_id;
  assign io_outputs_2_ar_validPipe_payload_len_1 = io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_len;
  assign io_outputs_2_ar_validPipe_payload_size_1 = io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_size;
  assign io_outputs_2_ar_validPipe_payload_burst_1 = io_axiOut_readOnly_decoder_1_io_outputs_2_ar_payload_burst;
  assign io_outputs_2_ar_validPipe_ready_1 = axi4ReadOnlyArbiter_5_io_inputs_1_ar_ready;
  assign io_axiOut_readOnly_decoder_1_io_outputs_2_r_payload_id = axi4ReadOnlyArbiter_5_io_inputs_1_r_payload_id[3:0];
  assign io_axiOut_readOnly_ar_ready_1 = io_axiOut_readOnly_decoder_1_io_input_ar_ready;
  assign io_axiOut_readOnly_r_valid_1 = io_axiOut_readOnly_decoder_1_io_input_r_valid;
  assign io_axiOut_readOnly_r_payload_data_1 = io_axiOut_readOnly_decoder_1_io_input_r_payload_data;
  assign io_axiOut_readOnly_r_payload_last_1 = io_axiOut_readOnly_decoder_1_io_input_r_payload_last;
  assign io_axiOut_readOnly_r_payload_id_1 = io_axiOut_readOnly_decoder_1_io_input_r_payload_id;
  assign io_axiOut_readOnly_r_payload_resp_1 = io_axiOut_readOnly_decoder_1_io_input_r_payload_resp;
  assign io_outputs_0_aw_validPipe_fire_1 = (io_outputs_0_aw_validPipe_valid_1 && io_outputs_0_aw_validPipe_ready_1);
  assign io_outputs_0_aw_validPipe_valid_1 = io_outputs_0_aw_rValid_1;
  assign io_outputs_0_aw_validPipe_payload_addr_1 = io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_addr;
  assign io_outputs_0_aw_validPipe_payload_id_1 = io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_id;
  assign io_outputs_0_aw_validPipe_payload_len_1 = io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_len;
  assign io_outputs_0_aw_validPipe_payload_size_1 = io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_size;
  assign io_outputs_0_aw_validPipe_payload_burst_1 = io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_payload_burst;
  assign io_outputs_0_aw_validPipe_ready_1 = axi4WriteOnlyArbiter_3_io_inputs_1_aw_ready;
  assign io_axiOut_writeOnly_decoder_1_io_outputs_0_b_payload_id = axi4WriteOnlyArbiter_3_io_inputs_1_b_payload_id[3:0];
  assign io_outputs_1_aw_validPipe_fire_1 = (io_outputs_1_aw_validPipe_valid_1 && io_outputs_1_aw_validPipe_ready_1);
  assign io_outputs_1_aw_validPipe_valid_1 = io_outputs_1_aw_rValid_1;
  assign io_outputs_1_aw_validPipe_payload_addr_1 = io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_addr;
  assign io_outputs_1_aw_validPipe_payload_id_1 = io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_id;
  assign io_outputs_1_aw_validPipe_payload_len_1 = io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_len;
  assign io_outputs_1_aw_validPipe_payload_size_1 = io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_size;
  assign io_outputs_1_aw_validPipe_payload_burst_1 = io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_payload_burst;
  assign io_outputs_1_aw_validPipe_ready_1 = axi4WriteOnlyArbiter_4_io_inputs_1_aw_ready;
  assign io_axiOut_writeOnly_decoder_1_io_outputs_1_b_payload_id = axi4WriteOnlyArbiter_4_io_inputs_1_b_payload_id[3:0];
  assign io_outputs_2_aw_validPipe_fire_1 = (io_outputs_2_aw_validPipe_valid_1 && io_outputs_2_aw_validPipe_ready_1);
  assign io_outputs_2_aw_validPipe_valid_1 = io_outputs_2_aw_rValid_1;
  assign io_outputs_2_aw_validPipe_payload_addr_1 = io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_addr;
  assign io_outputs_2_aw_validPipe_payload_id_1 = io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_id;
  assign io_outputs_2_aw_validPipe_payload_len_1 = io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_len;
  assign io_outputs_2_aw_validPipe_payload_size_1 = io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_size;
  assign io_outputs_2_aw_validPipe_payload_burst_1 = io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_payload_burst;
  assign io_outputs_2_aw_validPipe_ready_1 = axi4WriteOnlyArbiter_5_io_inputs_1_aw_ready;
  assign io_axiOut_writeOnly_decoder_1_io_outputs_2_b_payload_id = axi4WriteOnlyArbiter_5_io_inputs_1_b_payload_id[3:0];
  assign io_axiOut_writeOnly_aw_ready_1 = io_axiOut_writeOnly_decoder_1_io_input_aw_ready;
  assign io_axiOut_writeOnly_w_ready_1 = io_axiOut_writeOnly_decoder_1_io_input_w_ready;
  assign io_axiOut_writeOnly_b_valid_1 = io_axiOut_writeOnly_decoder_1_io_input_b_valid;
  assign io_axiOut_writeOnly_b_payload_id_1 = io_axiOut_writeOnly_decoder_1_io_input_b_payload_id;
  assign io_axiOut_writeOnly_b_payload_resp_1 = io_axiOut_writeOnly_decoder_1_io_input_b_payload_resp;
  assign io_outputs_0_ar_validPipe_fire_2 = (io_outputs_0_ar_validPipe_valid_2 && io_outputs_0_ar_validPipe_ready_2);
  assign io_outputs_0_ar_validPipe_valid_2 = io_outputs_0_ar_rValid_2;
  assign io_outputs_0_ar_validPipe_payload_addr_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_addr;
  assign io_outputs_0_ar_validPipe_payload_id_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_id;
  assign io_outputs_0_ar_validPipe_payload_len_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_len;
  assign io_outputs_0_ar_validPipe_payload_size_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_size;
  assign io_outputs_0_ar_validPipe_payload_burst_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_burst;
  assign io_outputs_0_ar_validPipe_payload_prot = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_payload_prot;
  assign io_outputs_0_ar_validPipe_ready_2 = axi4ReadOnlyArbiter_3_io_inputs_2_ar_ready;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_r_payload_id = axi4ReadOnlyArbiter_3_io_inputs_2_r_payload_id[2:0];
  assign io_outputs_1_ar_validPipe_fire_2 = (io_outputs_1_ar_validPipe_valid_2 && io_outputs_1_ar_validPipe_ready_2);
  assign io_outputs_1_ar_validPipe_valid_2 = io_outputs_1_ar_rValid_2;
  assign io_outputs_1_ar_validPipe_payload_addr_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_addr;
  assign io_outputs_1_ar_validPipe_payload_id_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_id;
  assign io_outputs_1_ar_validPipe_payload_len_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_len;
  assign io_outputs_1_ar_validPipe_payload_size_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_size;
  assign io_outputs_1_ar_validPipe_payload_burst_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_burst;
  assign io_outputs_1_ar_validPipe_payload_prot = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_payload_prot;
  assign io_outputs_1_ar_validPipe_ready_2 = axi4ReadOnlyArbiter_4_io_inputs_2_ar_ready;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_r_payload_id = axi4ReadOnlyArbiter_4_io_inputs_2_r_payload_id[2:0];
  assign io_outputs_2_ar_validPipe_fire_2 = (io_outputs_2_ar_validPipe_valid_2 && io_outputs_2_ar_validPipe_ready_2);
  assign io_outputs_2_ar_validPipe_valid_2 = io_outputs_2_ar_rValid_2;
  assign io_outputs_2_ar_validPipe_payload_addr_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_addr;
  assign io_outputs_2_ar_validPipe_payload_id_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_id;
  assign io_outputs_2_ar_validPipe_payload_len_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_len;
  assign io_outputs_2_ar_validPipe_payload_size_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_size;
  assign io_outputs_2_ar_validPipe_payload_burst_2 = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_burst;
  assign io_outputs_2_ar_validPipe_payload_prot = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_payload_prot;
  assign io_outputs_2_ar_validPipe_ready_2 = axi4ReadOnlyArbiter_5_io_inputs_2_ar_ready;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_r_payload_id = axi4ReadOnlyArbiter_5_io_inputs_2_r_payload_id[2:0];
  assign DataCachePlugin_setup_dcacheMaster_readOnly_ar_ready = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_ar_ready;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_r_valid = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_valid;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_data = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_data;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_last = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_last;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_id = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_id;
  assign DataCachePlugin_setup_dcacheMaster_readOnly_r_payload_resp = DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_input_r_payload_resp;
  assign io_outputs_0_aw_validPipe_fire_2 = (io_outputs_0_aw_validPipe_valid_2 && io_outputs_0_aw_validPipe_ready_2);
  assign io_outputs_0_aw_validPipe_valid_2 = io_outputs_0_aw_rValid_2;
  assign io_outputs_0_aw_validPipe_payload_addr_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  assign io_outputs_0_aw_validPipe_payload_id_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_id;
  assign io_outputs_0_aw_validPipe_payload_len_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_len;
  assign io_outputs_0_aw_validPipe_payload_size_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_size;
  assign io_outputs_0_aw_validPipe_payload_burst_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  assign io_outputs_0_aw_validPipe_payload_prot = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_payload_prot;
  assign io_outputs_0_aw_validPipe_ready_2 = axi4WriteOnlyArbiter_3_io_inputs_2_aw_ready;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_b_payload_id = axi4WriteOnlyArbiter_3_io_inputs_2_b_payload_id[2:0];
  assign io_outputs_1_aw_validPipe_fire_2 = (io_outputs_1_aw_validPipe_valid_2 && io_outputs_1_aw_validPipe_ready_2);
  assign io_outputs_1_aw_validPipe_valid_2 = io_outputs_1_aw_rValid_2;
  assign io_outputs_1_aw_validPipe_payload_addr_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_addr;
  assign io_outputs_1_aw_validPipe_payload_id_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_id;
  assign io_outputs_1_aw_validPipe_payload_len_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_len;
  assign io_outputs_1_aw_validPipe_payload_size_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_size;
  assign io_outputs_1_aw_validPipe_payload_burst_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_burst;
  assign io_outputs_1_aw_validPipe_payload_prot = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_payload_prot;
  assign io_outputs_1_aw_validPipe_ready_2 = axi4WriteOnlyArbiter_4_io_inputs_2_aw_ready;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_b_payload_id = axi4WriteOnlyArbiter_4_io_inputs_2_b_payload_id[2:0];
  assign io_outputs_2_aw_validPipe_fire_2 = (io_outputs_2_aw_validPipe_valid_2 && io_outputs_2_aw_validPipe_ready_2);
  assign io_outputs_2_aw_validPipe_valid_2 = io_outputs_2_aw_rValid_2;
  assign io_outputs_2_aw_validPipe_payload_addr_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_addr;
  assign io_outputs_2_aw_validPipe_payload_id_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_id;
  assign io_outputs_2_aw_validPipe_payload_len_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_len;
  assign io_outputs_2_aw_validPipe_payload_size_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_size;
  assign io_outputs_2_aw_validPipe_payload_burst_2 = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_burst;
  assign io_outputs_2_aw_validPipe_payload_prot = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_payload_prot;
  assign io_outputs_2_aw_validPipe_ready_2 = axi4WriteOnlyArbiter_5_io_inputs_2_aw_ready;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_b_payload_id = axi4WriteOnlyArbiter_5_io_inputs_2_b_payload_id[2:0];
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_aw_ready = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_aw_ready;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_w_ready = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_w_ready;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_b_valid = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_valid;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_b_payload_id = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_payload_id;
  assign DataCachePlugin_setup_dcacheMaster_writeOnly_b_payload_resp = DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_input_b_payload_resp;
  assign io_outputs_0_ar_validPipe_fire_3 = (io_outputs_0_ar_validPipe_valid_3 && io_outputs_0_ar_validPipe_ready_3);
  assign io_outputs_0_ar_validPipe_valid_3 = io_outputs_0_ar_rValid_3;
  assign io_outputs_0_ar_validPipe_payload_addr_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_addr;
  assign io_outputs_0_ar_validPipe_payload_id_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_id;
  assign io_outputs_0_ar_validPipe_payload_len_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_len;
  assign io_outputs_0_ar_validPipe_payload_size_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_size;
  assign io_outputs_0_ar_validPipe_payload_burst_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_payload_burst;
  assign io_outputs_0_ar_validPipe_ready_3 = axi4ReadOnlyArbiter_3_io_inputs_3_ar_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_r_payload_id = axi4ReadOnlyArbiter_3_io_inputs_3_r_payload_id[3:0];
  assign io_outputs_1_ar_validPipe_fire_3 = (io_outputs_1_ar_validPipe_valid_3 && io_outputs_1_ar_validPipe_ready_3);
  assign io_outputs_1_ar_validPipe_valid_3 = io_outputs_1_ar_rValid_3;
  assign io_outputs_1_ar_validPipe_payload_addr_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_addr;
  assign io_outputs_1_ar_validPipe_payload_id_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_id;
  assign io_outputs_1_ar_validPipe_payload_len_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_len;
  assign io_outputs_1_ar_validPipe_payload_size_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_size;
  assign io_outputs_1_ar_validPipe_payload_burst_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_payload_burst;
  assign io_outputs_1_ar_validPipe_ready_3 = axi4ReadOnlyArbiter_4_io_inputs_3_ar_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_r_payload_id = axi4ReadOnlyArbiter_4_io_inputs_3_r_payload_id[3:0];
  assign io_outputs_2_ar_validPipe_fire_3 = (io_outputs_2_ar_validPipe_valid_3 && io_outputs_2_ar_validPipe_ready_3);
  assign io_outputs_2_ar_validPipe_valid_3 = io_outputs_2_ar_rValid_3;
  assign io_outputs_2_ar_validPipe_payload_addr_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_addr;
  assign io_outputs_2_ar_validPipe_payload_id_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_id;
  assign io_outputs_2_ar_validPipe_payload_len_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_len;
  assign io_outputs_2_ar_validPipe_payload_size_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_size;
  assign io_outputs_2_ar_validPipe_payload_burst_3 = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_payload_burst;
  assign io_outputs_2_ar_validPipe_ready_3 = axi4ReadOnlyArbiter_5_io_inputs_3_ar_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_r_payload_id = axi4ReadOnlyArbiter_5_io_inputs_3_r_payload_id[3:0];
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_ar_ready = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_ar_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_r_valid = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_valid;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_data = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_data;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_last = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_last;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_id = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_id;
  assign CoreMemSysPlugin_logic_roMasters_0_readOnly_r_payload_resp = CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_input_r_payload_resp;
  assign io_outputs_0_aw_validPipe_fire_3 = (io_outputs_0_aw_validPipe_valid_3 && io_outputs_0_aw_validPipe_ready_3);
  assign io_outputs_0_aw_validPipe_valid_3 = io_outputs_0_aw_rValid_3;
  assign io_outputs_0_aw_validPipe_payload_addr_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  assign io_outputs_0_aw_validPipe_payload_id_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_id;
  assign io_outputs_0_aw_validPipe_payload_len_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_len;
  assign io_outputs_0_aw_validPipe_payload_size_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_size;
  assign io_outputs_0_aw_validPipe_payload_burst_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  assign io_outputs_0_aw_validPipe_ready_3 = axi4WriteOnlyArbiter_3_io_inputs_3_aw_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_b_payload_id = axi4WriteOnlyArbiter_3_io_inputs_3_b_payload_id[3:0];
  assign io_outputs_1_aw_validPipe_fire_3 = (io_outputs_1_aw_validPipe_valid_3 && io_outputs_1_aw_validPipe_ready_3);
  assign io_outputs_1_aw_validPipe_valid_3 = io_outputs_1_aw_rValid_3;
  assign io_outputs_1_aw_validPipe_payload_addr_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_addr;
  assign io_outputs_1_aw_validPipe_payload_id_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_id;
  assign io_outputs_1_aw_validPipe_payload_len_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_len;
  assign io_outputs_1_aw_validPipe_payload_size_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_size;
  assign io_outputs_1_aw_validPipe_payload_burst_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_payload_burst;
  assign io_outputs_1_aw_validPipe_ready_3 = axi4WriteOnlyArbiter_4_io_inputs_3_aw_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_b_payload_id = axi4WriteOnlyArbiter_4_io_inputs_3_b_payload_id[3:0];
  assign io_outputs_2_aw_validPipe_fire_3 = (io_outputs_2_aw_validPipe_valid_3 && io_outputs_2_aw_validPipe_ready_3);
  assign io_outputs_2_aw_validPipe_valid_3 = io_outputs_2_aw_rValid_3;
  assign io_outputs_2_aw_validPipe_payload_addr_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_addr;
  assign io_outputs_2_aw_validPipe_payload_id_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_id;
  assign io_outputs_2_aw_validPipe_payload_len_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_len;
  assign io_outputs_2_aw_validPipe_payload_size_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_size;
  assign io_outputs_2_aw_validPipe_payload_burst_3 = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_payload_burst;
  assign io_outputs_2_aw_validPipe_ready_3 = axi4WriteOnlyArbiter_5_io_inputs_3_aw_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_b_payload_id = axi4WriteOnlyArbiter_5_io_inputs_3_b_payload_id[3:0];
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_aw_ready = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_aw_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_w_ready = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_w_ready;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_valid = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_valid;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_payload_id = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_payload_id;
  assign CoreMemSysPlugin_logic_roMasters_0_writeOnly_b_payload_resp = CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_input_b_payload_resp;
  assign axi4ReadOnlyArbiter_3_io_inputs_0_ar_payload_id = {1'd0, io_outputs_0_ar_validPipe_payload_id};
  assign axi4ReadOnlyArbiter_3_io_inputs_1_ar_payload_id = {1'd0, io_outputs_0_ar_validPipe_payload_id_1};
  assign axi4ReadOnlyArbiter_3_io_inputs_2_ar_payload_id = {2'd0, io_outputs_0_ar_validPipe_payload_id_2};
  assign axi4ReadOnlyArbiter_3_io_inputs_3_ar_payload_id = {1'd0, io_outputs_0_ar_validPipe_payload_id_3};
  assign axi4WriteOnlyArbiter_3_io_inputs_0_aw_payload_id = {1'd0, io_outputs_0_aw_validPipe_payload_id};
  assign axi4WriteOnlyArbiter_3_io_inputs_1_aw_payload_id = {1'd0, io_outputs_0_aw_validPipe_payload_id_1};
  assign axi4WriteOnlyArbiter_3_io_inputs_2_aw_payload_id = {2'd0, io_outputs_0_aw_validPipe_payload_id_2};
  assign axi4WriteOnlyArbiter_3_io_inputs_3_aw_payload_id = {1'd0, io_outputs_0_aw_validPipe_payload_id_3};
  assign axi4ReadOnlyArbiter_4_io_inputs_0_ar_payload_id = {1'd0, io_outputs_1_ar_validPipe_payload_id};
  assign axi4ReadOnlyArbiter_4_io_inputs_1_ar_payload_id = {1'd0, io_outputs_1_ar_validPipe_payload_id_1};
  assign axi4ReadOnlyArbiter_4_io_inputs_2_ar_payload_id = {2'd0, io_outputs_1_ar_validPipe_payload_id_2};
  assign axi4ReadOnlyArbiter_4_io_inputs_3_ar_payload_id = {1'd0, io_outputs_1_ar_validPipe_payload_id_3};
  assign axi4WriteOnlyArbiter_4_io_inputs_0_aw_payload_id = {1'd0, io_outputs_1_aw_validPipe_payload_id};
  assign axi4WriteOnlyArbiter_4_io_inputs_1_aw_payload_id = {1'd0, io_outputs_1_aw_validPipe_payload_id_1};
  assign axi4WriteOnlyArbiter_4_io_inputs_2_aw_payload_id = {2'd0, io_outputs_1_aw_validPipe_payload_id_2};
  assign axi4WriteOnlyArbiter_4_io_inputs_3_aw_payload_id = {1'd0, io_outputs_1_aw_validPipe_payload_id_3};
  assign axi4ReadOnlyArbiter_5_io_inputs_0_ar_payload_id = {1'd0, io_outputs_2_ar_validPipe_payload_id};
  assign axi4ReadOnlyArbiter_5_io_inputs_1_ar_payload_id = {1'd0, io_outputs_2_ar_validPipe_payload_id_1};
  assign axi4ReadOnlyArbiter_5_io_inputs_2_ar_payload_id = {2'd0, io_outputs_2_ar_validPipe_payload_id_2};
  assign axi4ReadOnlyArbiter_5_io_inputs_3_ar_payload_id = {1'd0, io_outputs_2_ar_validPipe_payload_id_3};
  assign axi4WriteOnlyArbiter_5_io_inputs_0_aw_payload_id = {1'd0, io_outputs_2_aw_validPipe_payload_id};
  assign axi4WriteOnlyArbiter_5_io_inputs_1_aw_payload_id = {1'd0, io_outputs_2_aw_validPipe_payload_id_1};
  assign axi4WriteOnlyArbiter_5_io_inputs_2_aw_payload_id = {2'd0, io_outputs_2_aw_validPipe_payload_id_2};
  assign axi4WriteOnlyArbiter_5_io_inputs_3_aw_payload_id = {1'd0, io_outputs_2_aw_validPipe_payload_id_3};
  assign io_dpy0 = DebugDisplayPlugin_hw_dpyController_io_dpy0_out;
  assign io_dpy1 = DebugDisplayPlugin_hw_dpyController_io_dpy1_out;
  assign _zz_when_CoreNSCSCC_l598 = io_switch_btn_buffercc_io_dataOut;
  assign when_CoreNSCSCC_l598 = (_zz_when_CoreNSCSCC_l598 && (! _zz_when_CoreNSCSCC_l598_1));
  assign io_leds = _zz_io_leds_1[15:0];
  always @(posedge clk) begin
    if(reset) begin
      FetchPipelinePlugin_dbg_cycles <= 16'h0;
      FetchPipelinePlugin_dbg_c <= 3'b000;
      CommitPlugin_commitStatsReg_committedThisCycle <= 1'b0;
      CommitPlugin_commitStatsReg_totalCommitted <= 32'h0;
      CommitPlugin_commitStatsReg_robFlushCount <= 32'h0;
      CommitPlugin_commitStatsReg_physRegRecycled <= 32'h0;
      CommitPlugin_commitStatsReg_commitOOB <= 1'b0;
      CommitPlugin_commitStatsReg_maxCommitPc <= 32'h0;
      CommitPlugin_maxCommitPcReg <= 32'h0;
      CommitPlugin_commitOOBReg <= 1'b0;
      _zz_when_Debug_l71 <= 8'h0;
      io_mem_read_cmd_rValid <= 1'b0;
      DataCachePlugin_setup_dcacheMaster_r_rValid <= 1'b0;
      io_mem_write_cmd_fork2_logic_linkEnable_0 <= 1'b1;
      io_mem_write_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      io_mem_toAxi4_awRaw_payload_first <= 1'b1;
      io_mem_toAxi4_awFiltred_rValid <= 1'b0;
      io_mem_toAxi4_w_rValid <= 1'b0;
      DataCachePlugin_setup_dcacheMaster_b_rValid <= 1'b0;
      BusyTablePlugin_early_setup_busyTableReg <= 64'h0;
      CheckpointManagerPlugin_logic_hasValidCheckpoint <= 1'b0;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_0 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_0;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_1 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_1;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_2 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_2;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_3 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_3;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_4 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_4;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_5 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_5;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_6 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_6;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_7 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_7;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_8 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_8;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_9 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_9;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_10 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_10;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_11 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_11;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_12 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_12;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_13 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_13;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_14 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_14;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_15 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_15;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_16 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_16;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_17 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_17;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_18 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_18;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_19 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_19;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_20 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_20;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_21 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_21;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_22 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_22;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_23 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_23;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_24 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_24;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_25 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_25;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_26 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_26;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_27 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_27;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_28 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_28;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_29 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_29;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_30 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_30;
      CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_31 <= CheckpointManagerPlugin_logic_initialRatCheckpoint_mapping_31;
      CheckpointManagerPlugin_logic_storedBtCheckpoint_busyBits <= CheckpointManagerPlugin_logic_initialBtCheckpoint_busyBits;
      CommitPlugin_logic_s1_s1_committedThisCycle <= 1'b0;
      CommitPlugin_logic_s1_s1_recycledThisCycle <= 1'b0;
      CommitPlugin_logic_s1_s1_flushedThisCycle <= 1'b0;
      CommitPlugin_logic_s1_s1_maxCommitPcThisCycle <= 32'h0;
      CommitPlugin_logic_s1_s1_anyCommitOOB <= 1'b0;
      CommitPlugin_logic_counter <= 32'h0;
      DebugDisplayPlugin_logic_displayArea_dpToggle <= 1'b0;
      s1_ReadRegs_valid <= 1'b0;
      s2_Execute_valid <= 1'b0;
      s3_Writeback_valid <= 1'b0;
      mul_s1_ReadRegs_valid <= 1'b0;
      mul_s2_Execute_valid <= 1'b0;
      mul_s3_Execute_valid <= 1'b0;
      mul_s4_Execute_valid <= 1'b0;
      mul_s5_Execute_valid <= 1'b0;
      mul_s6_Execute_valid <= 1'b0;
      mul_s7_Writeback_valid <= 1'b0;
      s1_Calc_valid <= 1'b0;
      s2_Select_valid <= 1'b0;
      s3_Result_valid <= 1'b0;
      s1_Rename_valid <= 1'b0;
      s2_RobAlloc_valid <= 1'b0;
      s3_Dispatch_valid <= 1'b0;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid <= 1'b0;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid_2 <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromFwd <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromDCache <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromMMIO <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromEarlyExc <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_data <= 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_hasFault <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_exceptionCode <= 8'bxxxxxxxx;
      LoadQueuePlugin_logic_loadQueue_sbQueryRspValid <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_registeredFlush_valid <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr <= 4'b0000;
      LoadQueuePlugin_logic_loadQueue_slots_0_valid <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_0_address <= 32'h0;
      LoadQueuePlugin_logic_loadQueue_slots_0_size <= MemAccessSize_W;
      LoadQueuePlugin_logic_loadQueue_slots_0_robPtr <= 4'b0000;
      LoadQueuePlugin_logic_loadQueue_slots_0_pdest <= 6'h0;
      LoadQueuePlugin_logic_loadQueue_slots_0_isIO <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_0_hasException <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_0_exceptionCode <= 8'h0;
      LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_0_isStalledByDependency <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_1_valid <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_1_address <= 32'h0;
      LoadQueuePlugin_logic_loadQueue_slots_1_size <= MemAccessSize_W;
      LoadQueuePlugin_logic_loadQueue_slots_1_robPtr <= 4'b0000;
      LoadQueuePlugin_logic_loadQueue_slots_1_pdest <= 6'h0;
      LoadQueuePlugin_logic_loadQueue_slots_1_isIO <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_1_hasException <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_1_exceptionCode <= 8'h0;
      LoadQueuePlugin_logic_loadQueue_slots_1_isWaitingForFwdRsp <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_1_isStalledByDependency <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_1_isReadyForDCache <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_1_isWaitingForRsp <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_2_valid <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_2_address <= 32'h0;
      LoadQueuePlugin_logic_loadQueue_slots_2_size <= MemAccessSize_W;
      LoadQueuePlugin_logic_loadQueue_slots_2_robPtr <= 4'b0000;
      LoadQueuePlugin_logic_loadQueue_slots_2_pdest <= 6'h0;
      LoadQueuePlugin_logic_loadQueue_slots_2_isIO <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_2_hasException <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_2_exceptionCode <= 8'h0;
      LoadQueuePlugin_logic_loadQueue_slots_2_isWaitingForFwdRsp <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_2_isStalledByDependency <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_2_isReadyForDCache <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_2_isWaitingForRsp <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_3_valid <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_3_address <= 32'h0;
      LoadQueuePlugin_logic_loadQueue_slots_3_size <= MemAccessSize_W;
      LoadQueuePlugin_logic_loadQueue_slots_3_robPtr <= 4'b0000;
      LoadQueuePlugin_logic_loadQueue_slots_3_pdest <= 6'h0;
      LoadQueuePlugin_logic_loadQueue_slots_3_isIO <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_3_hasException <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_3_exceptionCode <= 8'h0;
      LoadQueuePlugin_logic_loadQueue_slots_3_isWaitingForFwdRsp <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_3_isStalledByDependency <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_3_isReadyForDCache <= 1'b0;
      LoadQueuePlugin_logic_loadQueue_slots_3_isWaitingForRsp <= 1'b0;
      PhysicalRegFilePlugin_logic_regFile_0 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_1 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_2 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_3 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_4 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_5 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_6 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_7 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_8 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_9 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_10 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_11 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_12 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_13 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_14 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_15 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_16 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_17 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_18 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_19 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_20 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_21 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_22 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_23 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_24 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_25 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_26 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_27 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_28 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_29 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_30 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_31 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_32 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_33 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_34 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_35 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_36 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_37 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_38 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_39 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_40 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_41 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_42 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_43 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_44 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_45 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_46 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_47 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_48 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_49 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_50 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_51 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_52 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_53 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_54 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_55 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_56 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_57 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_58 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_59 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_60 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_61 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_62 <= 32'h0;
      PhysicalRegFilePlugin_logic_regFile_63 <= 32'h0;
      StoreBufferPlugin_logic_slots_0_isFlush <= 1'b0;
      StoreBufferPlugin_logic_slots_0_addr <= 32'h0;
      StoreBufferPlugin_logic_slots_0_data <= 32'h0;
      StoreBufferPlugin_logic_slots_0_be <= 4'b0000;
      StoreBufferPlugin_logic_slots_0_robPtr <= 4'b0000;
      StoreBufferPlugin_logic_slots_0_accessSize <= MemAccessSize_W;
      StoreBufferPlugin_logic_slots_0_isIO <= 1'b0;
      StoreBufferPlugin_logic_slots_0_valid <= 1'b0;
      StoreBufferPlugin_logic_slots_0_hasEarlyException <= 1'b0;
      StoreBufferPlugin_logic_slots_0_earlyExceptionCode <= 8'h0;
      StoreBufferPlugin_logic_slots_0_isCommitted <= 1'b0;
      StoreBufferPlugin_logic_slots_0_sentCmd <= 1'b0;
      StoreBufferPlugin_logic_slots_0_waitRsp <= 1'b0;
      StoreBufferPlugin_logic_slots_0_isWaitingForRefill <= 1'b0;
      StoreBufferPlugin_logic_slots_0_isWaitingForWb <= 1'b0;
      StoreBufferPlugin_logic_slots_0_refillSlotToWatch <= 8'h0;
      StoreBufferPlugin_logic_slots_1_isFlush <= 1'b0;
      StoreBufferPlugin_logic_slots_1_addr <= 32'h0;
      StoreBufferPlugin_logic_slots_1_data <= 32'h0;
      StoreBufferPlugin_logic_slots_1_be <= 4'b0000;
      StoreBufferPlugin_logic_slots_1_robPtr <= 4'b0000;
      StoreBufferPlugin_logic_slots_1_accessSize <= MemAccessSize_W;
      StoreBufferPlugin_logic_slots_1_isIO <= 1'b0;
      StoreBufferPlugin_logic_slots_1_valid <= 1'b0;
      StoreBufferPlugin_logic_slots_1_hasEarlyException <= 1'b0;
      StoreBufferPlugin_logic_slots_1_earlyExceptionCode <= 8'h0;
      StoreBufferPlugin_logic_slots_1_isCommitted <= 1'b0;
      StoreBufferPlugin_logic_slots_1_sentCmd <= 1'b0;
      StoreBufferPlugin_logic_slots_1_waitRsp <= 1'b0;
      StoreBufferPlugin_logic_slots_1_isWaitingForRefill <= 1'b0;
      StoreBufferPlugin_logic_slots_1_isWaitingForWb <= 1'b0;
      StoreBufferPlugin_logic_slots_1_refillSlotToWatch <= 8'h0;
      StoreBufferPlugin_logic_slots_2_isFlush <= 1'b0;
      StoreBufferPlugin_logic_slots_2_addr <= 32'h0;
      StoreBufferPlugin_logic_slots_2_data <= 32'h0;
      StoreBufferPlugin_logic_slots_2_be <= 4'b0000;
      StoreBufferPlugin_logic_slots_2_robPtr <= 4'b0000;
      StoreBufferPlugin_logic_slots_2_accessSize <= MemAccessSize_W;
      StoreBufferPlugin_logic_slots_2_isIO <= 1'b0;
      StoreBufferPlugin_logic_slots_2_valid <= 1'b0;
      StoreBufferPlugin_logic_slots_2_hasEarlyException <= 1'b0;
      StoreBufferPlugin_logic_slots_2_earlyExceptionCode <= 8'h0;
      StoreBufferPlugin_logic_slots_2_isCommitted <= 1'b0;
      StoreBufferPlugin_logic_slots_2_sentCmd <= 1'b0;
      StoreBufferPlugin_logic_slots_2_waitRsp <= 1'b0;
      StoreBufferPlugin_logic_slots_2_isWaitingForRefill <= 1'b0;
      StoreBufferPlugin_logic_slots_2_isWaitingForWb <= 1'b0;
      StoreBufferPlugin_logic_slots_2_refillSlotToWatch <= 8'h0;
      StoreBufferPlugin_logic_slots_3_isFlush <= 1'b0;
      StoreBufferPlugin_logic_slots_3_addr <= 32'h0;
      StoreBufferPlugin_logic_slots_3_data <= 32'h0;
      StoreBufferPlugin_logic_slots_3_be <= 4'b0000;
      StoreBufferPlugin_logic_slots_3_robPtr <= 4'b0000;
      StoreBufferPlugin_logic_slots_3_accessSize <= MemAccessSize_W;
      StoreBufferPlugin_logic_slots_3_isIO <= 1'b0;
      StoreBufferPlugin_logic_slots_3_valid <= 1'b0;
      StoreBufferPlugin_logic_slots_3_hasEarlyException <= 1'b0;
      StoreBufferPlugin_logic_slots_3_earlyExceptionCode <= 8'h0;
      StoreBufferPlugin_logic_slots_3_isCommitted <= 1'b0;
      StoreBufferPlugin_logic_slots_3_sentCmd <= 1'b0;
      StoreBufferPlugin_logic_slots_3_waitRsp <= 1'b0;
      StoreBufferPlugin_logic_slots_3_isWaitingForRefill <= 1'b0;
      StoreBufferPlugin_logic_slots_3_isWaitingForWb <= 1'b0;
      StoreBufferPlugin_logic_slots_3_refillSlotToWatch <= 8'h0;
      StoreBufferPlugin_logic_registeredFlush_valid <= 1'b0;
      StoreBufferPlugin_logic_registeredFlush_targetRobPtr <= 4'b0000;
      StoreBufferPlugin_logic_registeredCommitUpdate_validMask <= 4'b0000;
      FetchPipelinePlugin_logic_retryIdCounter_value <= 2'b01;
      FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value <= 3'b000;
      FetchPipelinePlugin_logic_isDrainingCacheRspReg <= 1'b0;
      FetchPipelinePlugin_logic_retryCmd_lock <= 1'b0;
      FetchPipelinePlugin_logic_retryCmd_pc <= 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      FetchPipelinePlugin_logic_retryCmd_id <= 2'bxx;
      FetchPipelinePlugin_logic_s1_logic_fetchPcReg <= 32'h80000000;
      FetchPipelinePlugin_logic_s1_logic_lastRetryIdReg <= 2'b00;
      s2_ICache_Access_valid <= 1'b0;
      s4_Predecode_valid <= 1'b0;
      _zz_DataCachePlugin_logic_load_ohHistory_1 <= 1'b0;
      _zz_DataCachePlugin_logic_load_ohHistory_2 <= 1'b0;
      ICachePlugin_logic_storage_valids_0_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_0_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_1_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_1_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_2_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_2_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_3_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_3_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_4_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_4_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_5_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_5_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_6_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_6_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_7_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_7_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_8_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_8_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_9_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_9_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_10_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_10_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_11_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_11_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_12_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_12_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_13_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_13_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_14_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_14_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_15_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_15_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_16_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_16_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_17_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_17_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_18_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_18_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_19_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_19_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_20_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_20_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_21_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_21_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_22_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_22_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_23_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_23_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_24_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_24_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_25_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_25_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_26_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_26_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_27_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_27_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_28_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_28_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_29_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_29_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_30_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_30_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_31_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_31_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_32_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_32_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_33_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_33_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_34_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_34_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_35_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_35_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_36_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_36_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_37_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_37_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_38_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_38_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_39_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_39_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_40_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_40_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_41_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_41_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_42_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_42_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_43_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_43_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_44_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_44_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_45_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_45_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_46_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_46_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_47_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_47_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_48_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_48_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_49_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_49_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_50_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_50_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_51_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_51_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_52_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_52_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_53_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_53_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_54_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_54_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_55_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_55_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_56_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_56_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_57_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_57_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_58_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_58_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_59_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_59_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_60_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_60_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_61_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_61_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_62_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_62_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_63_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_63_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_64_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_64_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_65_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_65_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_66_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_66_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_67_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_67_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_68_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_68_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_69_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_69_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_70_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_70_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_71_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_71_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_72_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_72_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_73_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_73_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_74_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_74_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_75_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_75_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_76_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_76_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_77_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_77_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_78_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_78_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_79_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_79_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_80_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_80_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_81_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_81_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_82_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_82_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_83_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_83_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_84_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_84_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_85_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_85_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_86_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_86_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_87_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_87_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_88_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_88_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_89_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_89_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_90_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_90_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_91_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_91_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_92_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_92_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_93_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_93_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_94_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_94_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_95_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_95_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_96_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_96_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_97_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_97_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_98_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_98_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_99_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_99_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_100_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_100_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_101_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_101_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_102_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_102_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_103_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_103_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_104_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_104_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_105_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_105_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_106_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_106_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_107_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_107_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_108_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_108_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_109_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_109_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_110_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_110_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_111_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_111_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_112_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_112_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_113_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_113_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_114_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_114_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_115_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_115_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_116_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_116_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_117_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_117_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_118_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_118_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_119_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_119_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_120_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_120_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_121_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_121_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_122_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_122_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_123_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_123_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_124_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_124_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_125_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_125_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_126_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_126_1 <= 1'b0;
      ICachePlugin_logic_storage_valids_127_0 <= 1'b0;
      ICachePlugin_logic_storage_valids_127_1 <= 1'b0;
      ICachePlugin_logic_refill_refillCounter_value <= 2'b00;
      ICachePlugin_logic_refill_fsm_stateReg <= ICachePlugin_logic_refill_fsm_BOOT;
      ICache_F2_HitCheck_valid <= 1'b0;
      BpuPipelinePlugin_logic_s2_predict_valid <= 1'b0;
      BpuPipelinePlugin_logic_u2_write_valid <= 1'b0;
      io_outputs_0_ar_rValid <= 1'b0;
      io_outputs_1_ar_rValid <= 1'b0;
      io_outputs_2_ar_rValid <= 1'b0;
      io_outputs_0_aw_rValid <= 1'b0;
      io_outputs_1_aw_rValid <= 1'b0;
      io_outputs_2_aw_rValid <= 1'b0;
      io_outputs_0_ar_rValid_1 <= 1'b0;
      io_outputs_1_ar_rValid_1 <= 1'b0;
      io_outputs_2_ar_rValid_1 <= 1'b0;
      io_outputs_0_aw_rValid_1 <= 1'b0;
      io_outputs_1_aw_rValid_1 <= 1'b0;
      io_outputs_2_aw_rValid_1 <= 1'b0;
      io_outputs_0_ar_rValid_2 <= 1'b0;
      io_outputs_1_ar_rValid_2 <= 1'b0;
      io_outputs_2_ar_rValid_2 <= 1'b0;
      io_outputs_0_aw_rValid_2 <= 1'b0;
      io_outputs_1_aw_rValid_2 <= 1'b0;
      io_outputs_2_aw_rValid_2 <= 1'b0;
      io_outputs_0_ar_rValid_3 <= 1'b0;
      io_outputs_1_ar_rValid_3 <= 1'b0;
      io_outputs_2_ar_rValid_3 <= 1'b0;
      io_outputs_0_aw_rValid_3 <= 1'b0;
      io_outputs_1_aw_rValid_3 <= 1'b0;
      io_outputs_2_aw_rValid_3 <= 1'b0;
      _zz_io_leds <= 1'b0;
    end else begin
      FetchPipelinePlugin_dbg_cycles <= (FetchPipelinePlugin_dbg_cycles + 16'h0001);
      FetchPipelinePlugin_dbg_c <= (FetchPipelinePlugin_dbg_c + 3'b001);
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // FetchPipelinePlugin2.scala:L135
        `else
          if(!1'b0) begin
            $display("NOTE(FetchPipelinePlugin2.scala:135):  [normal] ------------ End of cycle 0x%x", FetchPipelinePlugin_dbg_cycles); // FetchPipelinePlugin2.scala:L135
          end
        `endif
      `endif
      if(DataCachePlugin_setup_cache_io_mem_read_cmd_ready) begin
        io_mem_read_cmd_rValid <= DataCachePlugin_setup_cache_io_mem_read_cmd_valid;
      end
      if(DataCachePlugin_setup_dcacheMaster_r_ready) begin
        DataCachePlugin_setup_dcacheMaster_r_rValid <= DataCachePlugin_setup_dcacheMaster_r_valid;
      end
      if(io_mem_toAxi4_awRaw_fire) begin
        io_mem_write_cmd_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(io_mem_toAxi4_wRaw_fire) begin
        io_mem_write_cmd_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(DataCachePlugin_setup_cache_io_mem_write_cmd_ready) begin
        io_mem_write_cmd_fork2_logic_linkEnable_0 <= 1'b1;
        io_mem_write_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(io_mem_toAxi4_awRaw_fire) begin
        io_mem_toAxi4_awRaw_payload_first <= io_mem_toAxi4_awRaw_payload_last;
      end
      if(io_mem_toAxi4_awFiltred_ready) begin
        io_mem_toAxi4_awFiltred_rValid <= io_mem_toAxi4_awFiltred_valid;
      end
      if(io_mem_toAxi4_w_ready) begin
        io_mem_toAxi4_w_rValid <= io_mem_toAxi4_w_valid;
      end
      if(DataCachePlugin_setup_dcacheMaster_b_ready) begin
        DataCachePlugin_setup_dcacheMaster_b_rValid <= DataCachePlugin_setup_dcacheMaster_b_valid;
      end
      if(oneShot_13_io_pulseOut) begin
        if(when_Debug_l71) begin
          _zz_when_Debug_l71 <= {7'd0, _zz_when_Debug_l71_1};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_1); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(oneShot_14_io_pulseOut) begin
        if(when_Debug_l71_1) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_2};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_2); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(oneShot_15_io_pulseOut) begin
        if(when_Debug_l71_2) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_3};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_3); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(oneShot_16_io_pulseOut) begin
        if(when_Debug_l71_3) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_4};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_4); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(oneShot_17_io_pulseOut) begin
        if(when_Debug_l71_4) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_5};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_5); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(CheckpointManagerPlugin_saveCheckpointTrigger) begin
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_0 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_0;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_1 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_1;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_2 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_2;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_3 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_3;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_4 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_4;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_5 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_5;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_6 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_6;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_7 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_7;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_8 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_8;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_9 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_9;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_10 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_10;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_11 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_11;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_12 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_12;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_13 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_13;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_14 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_14;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_15 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_15;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_16 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_16;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_17 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_17;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_18 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_18;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_19 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_19;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_20 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_20;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_21 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_21;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_22 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_22;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_23 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_23;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_24 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_24;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_25 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_25;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_26 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_26;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_27 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_27;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_28 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_28;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_29 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_29;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_30 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_30;
        CheckpointManagerPlugin_logic_storedRatCheckpoint_mapping_31 <= RenameMapTablePlugin_early_setup_rat_io_currentState_mapping_31;
        CheckpointManagerPlugin_logic_storedBtCheckpoint_busyBits <= BusyTablePlugin_early_setup_busyTableReg;
        CheckpointManagerPlugin_logic_hasValidCheckpoint <= 1'b1;
      end
      if(when_CommitPlugin_l203) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // CommitPlugin.scala:L208
          `else
            if(!1'b0) begin
              $display("NOTE(CommitPlugin.scala:208):  [COMMIT] BPU UPDATE: pc=0x%x, isTaken=%x, target=0x%x", BpuPipelinePlugin_updatePortIn_payload_pc, BpuPipelinePlugin_updatePortIn_payload_isTaken, BpuPipelinePlugin_updatePortIn_payload_target); // CommitPlugin.scala:L208
            end
          `endif
        `endif
      end else begin
        if(ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isBranchOrJump) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // CommitPlugin.scala:L211
            `else
              if(!1'b0) begin
                $display("NOTE(CommitPlugin.scala:211):  [COMMIT] BPU Not upated because enable=%x headSlot.canCommit=%x headIsBranch=%x", CommitPlugin_commitEnableExt, ROBPlugin_robComponent_io_commit_0_canCommit, ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_isBranchOrJump); // CommitPlugin.scala:L211
              end
            `endif
          `endif
        end
      end
      if(when_CommitPlugin_l216) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // CommitPlugin.scala:L223
          `else
            if(!1'b0) begin
              $display("NOTE(CommitPlugin.scala:223):  CHECKPOINT: Save checkpoint triggered on successful commit."); // CommitPlugin.scala:L223
            end
          `endif
        `endif
      end
      if(when_CommitPlugin_l227) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // CommitPlugin.scala:L244
          `else
            if(!1'b0) begin
              $display("NOTE(CommitPlugin.scala:244):  [notice] [33mBRANCH MISPREDICT: Vetoing commit of robPtr=%x, PC=0x%x and flushing pipeline. Redirecting to 0x%x.[0m", ROBPlugin_robComponent_io_commit_0_entry_payload_uop_robPtr, ROBPlugin_robComponent_io_commit_0_entry_payload_uop_decoded_pc, ROBPlugin_robComponent_io_commit_0_entry_status_result); // CommitPlugin.scala:L244
            end
          `endif
        `endif
      end
      CommitPlugin_logic_s1_s1_committedThisCycle <= CommitPlugin_logic_s0_committedThisCycle_comb;
      CommitPlugin_logic_s1_s1_recycledThisCycle <= CommitPlugin_logic_s0_recycledThisCycle_comb;
      CommitPlugin_logic_s1_s1_flushedThisCycle <= CommitPlugin_logic_s0_flushedThisCycle_comb;
      CommitPlugin_logic_s1_s1_maxCommitPcThisCycle <= CommitPlugin_logic_s0_maxCommitPcThisCycle;
      CommitPlugin_logic_s1_s1_anyCommitOOB <= CommitPlugin_logic_s0_anyCommitOOB;
      if(when_CommitPlugin_l317) begin
        CommitPlugin_maxCommitPcReg <= CommitPlugin_logic_s1_s1_maxCommitPcThisCycle;
      end
      if(CommitPlugin_logic_s1_s1_anyCommitOOB) begin
        CommitPlugin_commitOOBReg <= 1'b1;
      end
      CommitPlugin_commitStatsReg_committedThisCycle <= CommitPlugin_logic_s1_s1_committedThisCycle;
      CommitPlugin_commitStatsReg_totalCommitted <= (CommitPlugin_commitStatsReg_totalCommitted + _zz_CommitPlugin_commitStatsReg_totalCommitted);
      CommitPlugin_commitStatsReg_physRegRecycled <= (CommitPlugin_commitStatsReg_physRegRecycled + _zz_CommitPlugin_commitStatsReg_physRegRecycled);
      CommitPlugin_commitStatsReg_robFlushCount <= (CommitPlugin_commitStatsReg_robFlushCount + _zz_CommitPlugin_commitStatsReg_robFlushCount);
      CommitPlugin_commitStatsReg_commitOOB <= CommitPlugin_commitOOBReg;
      CommitPlugin_commitStatsReg_maxCommitPc <= CommitPlugin_maxCommitPcReg;
      if(oneShot_18_io_pulseOut) begin
        if(when_Debug_l71_5) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_6};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_6); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(oneShot_19_io_pulseOut) begin
        _zz_when_Debug_l71 <= 8'he3;
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // Debug.scala:L77
          `else
            if(!1'b0) begin
              $display("NOTE(Debug.scala:77):  [DbgSvc] Set value to 0x%x", _zz_26); // Debug.scala:L77
            end
          `endif
        `endif
      end
      CommitPlugin_logic_counter <= (CommitPlugin_logic_counter + 32'h00000001);
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // CommitPlugin.scala:L349
        `else
          if(!1'b0) begin
            $display("NOTE(CommitPlugin.scala:349):  [COMMIT] Cycle %x Log: Stats=CommitStats(committedThisCycle=%x, totalCommitted=%x, robFlushCount=%x, physRegRecycled=%x, commitOOB=%x, maxCommitPc=0x%x)\n  Slot Details: \n    Slot: (valid=%x, canCommit=%x, doCommit=%x, robPtr=%x, oldPhysDest=%x, allocatesPhysDest=%x) commitAck=%x commitPc=0x%x", CommitPlugin_logic_counter, CommitPlugin_commitStatsReg_committedThisCycle, CommitPlugin_commitStatsReg_totalCommitted, CommitPlugin_commitStatsReg_robFlushCount, CommitPlugin_commitStatsReg_physRegRecycled, CommitPlugin_commitStatsReg_commitOOB, CommitPlugin_commitStatsReg_maxCommitPc, CommitPlugin_logic_s0_commitSlotLogs_0_valid, CommitPlugin_logic_s0_commitSlotLogs_0_canCommit, CommitPlugin_logic_s0_commitSlotLogs_0_doCommit, CommitPlugin_logic_s0_commitSlotLogs_0_robPtr, CommitPlugin_logic_s0_commitSlotLogs_0_oldPhysDest, CommitPlugin_logic_s0_commitSlotLogs_0_allocatesPhysDest, CommitPlugin_logic_s0_commitAckMasks_0, CommitPlugin_logic_s0_commitPcs_0); // CommitPlugin.scala:L349
          end
        `endif
      `endif
      if(when_DecodePlugin_l117) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // DecodePlugin.scala:L118
          `else
            if(!1'b0) begin
              $display("NOTE(DecodePlugin.scala:118):  DecodePlugin (s0_decode): Firing. Output DecodedUops=DecodedUop @ pc=%x (%x)\n  Core Info:   uopCode=%s  exeUnit=%s  isa=%s\n  Operands:\n    dest=ArchRegOperand: idx=%xrtype=%sisGPR=%xisFPR=%xisCSR=%x writeEn=%x\n    src1=ArchRegOperand: idx=%xrtype=%sisGPR=%xisFPR=%xisCSR=%x use=%x\n    src2=ArchRegOperand: idx=%xrtype=%sisGPR=%xisFPR=%xisCSR=%x use=%x\n use=\n    imm=%x (usage=%s)\n  Control Flags:\n    ALU: AluCtrlFlags: isSub=%x isAdd=%x isSigned=%x logicOp=%s\n    Shift: ShiftCtrlFlags: isRight=%x isArithmetic=%x isRotate=%x isDoubleWord=%x\n    MulDiv: MulDivCtrlFlags: isDiv=%x isSigned=%x isWordOp=%x\n    Mem: MemCtrlFlags: size=%s isSignedLoad=%x isStore=%x isLoadLinked=%x isStoreCond=%x atomicOp=%x isFence=%x fenceMode=%x isCacheOp=%x cacheOpType=%x isPrefetch=%x\n    Branch: BranchCtrlFlags: condition=%s isJump=%x isLink=%x linkReg=ArchRegOperand: idx=%xrtype=%sisGPR=%xisFPR=%xisCSR=%x isIndirect=%x laCfIdx=%x\n    FPU: FpuCtrlFlags: opType=%x fpSizeSrc1=%s fpSizeSrc2=%s fpSizeDest=%s roundingMode=%x isIntegerDest=%x isSignedCvt=%x fmaNegSrc1=%x fcmpCond=%x\n    CSR: CsrCtrlFlags: csrAddr=%x isWrite=%x isRead=%x isExchange=%x useUimmAsSrc=%x\n    System: SystemCtrlFlags: sysCode=%x isExceptionReturn=%x isTlbOp=%x tlbOpType=%x\n  Status:\n    decodeEx=%s hasEx=%x\n    isMicrocode=%x entry=%x\n    isSerializing=%x isBranchOrJump=%x branchPrediction=BranchPredictionInfo: isTaken=%x target=%x wasPredicted=%x", DecodePlugin_logic_decodedUopsOutputVec_0_pc, DecodePlugin_logic_decodedUopsOutputVec_0_isValid, DecodePlugin_logic_decodedUopsOutputVec_0_uopCode_string, DecodePlugin_logic_decodedUopsOutputVec_0_exeUnit_string, DecodePlugin_logic_decodedUopsOutputVec_0_isa_string, DecodePlugin_logic_decodedUopsOutputVec_0_archDest_idx, DecodePlugin_logic_decodedUopsOutputVec_0_archDest_rtype_string, _zz_27, _zz_28, _zz_29, DecodePlugin_logic_decodedUopsOutputVec_0_writeArchDestEn, DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_idx, DecodePlugin_logic_decodedUopsOutputVec_0_archSrc1_rtype_string, _zz_30, _zz_31, _zz_32, DecodePlugin_logic_decodedUopsOutputVec_0_useArchSrc1, DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_idx, DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype_string, _zz_33, _zz_34, _zz_35, DecodePlugin_logic_decodedUopsOutputVec_0_useArchSrc2, DecodePlugin_logic_decodedUopsOutputVec_0_imm, DecodePlugin_logic_decodedUopsOutputVec_0_immUsage_string, DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isSub, DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isAdd, DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_isSigned, DecodePlugin_logic_decodedUopsOutputVec_0_aluCtrl_logicOp_string, DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isRight, DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isArithmetic, DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isRotate, DecodePlugin_logic_decodedUopsOutputVec_0_shiftCtrl_isDoubleWord, DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isDiv, DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isSigned, DecodePlugin_logic_decodedUopsOutputVec_0_mulDivCtrl_isWordOp, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_size_string, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isSignedLoad, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isStore, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isLoadLinked, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isStoreCond, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_atomicOp, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isFence, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_fenceMode, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isCacheOp, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_cacheOpType, DecodePlugin_logic_decodedUopsOutputVec_0_memCtrl_isPrefetch, DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_condition_string, DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isJump, DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isLink, DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_idx, DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_linkReg_rtype_string, _zz_36, _zz_37, _zz_38, DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_isIndirect, DecodePlugin_logic_decodedUopsOutputVec_0_branchCtrl_laCfIdx, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_opType, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc1_string, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeSrc2_string, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fpSizeDest_string, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_roundingMode, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_isIntegerDest, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_isSignedCvt, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fmaNegSrc1, DecodePlugin_logic_decodedUopsOutputVec_0_fpuCtrl_fcmpCond, DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_csrAddr, DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isWrite, DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isRead, DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_isExchange, DecodePlugin_logic_decodedUopsOutputVec_0_csrCtrl_useUimmAsSrc, DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_sysCode, DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_isExceptionReturn, DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_isTlbOp, DecodePlugin_logic_decodedUopsOutputVec_0_sysCtrl_tlbOpType, DecodePlugin_logic_decodedUopsOutputVec_0_decodeExceptionCode_string, DecodePlugin_logic_decodedUopsOutputVec_0_hasDecodeException, DecodePlugin_logic_decodedUopsOutputVec_0_isMicrocode, DecodePlugin_logic_decodedUopsOutputVec_0_microcodeEntry, DecodePlugin_logic_decodedUopsOutputVec_0_isSerializing, DecodePlugin_logic_decodedUopsOutputVec_0_isBranchOrJump, DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_isTaken, DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_target, DecodePlugin_logic_decodedUopsOutputVec_0_branchPrediction_wasPredicted); // DecodePlugin.scala:L118
            end
          `endif
        `endif
      end
      if(when_RenamePlugin_l83) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // RenamePlugin.scala:L84
          `else
            if(!1'b0) begin
              $display("NOTE(RenamePlugin.scala:84):  [notice] [33mS2: Failed to allocate physical registers for uops: DecodedUop @ pc=%x (%x)\n  Core Info:   uopCode=%s  exeUnit=%s  isa=%s\n  Operands:\n    dest=ArchRegOperand: idx=%xrtype=%sisGPR=%xisFPR=%xisCSR=%x writeEn=%x\n    src1=ArchRegOperand: idx=%xrtype=%sisGPR=%xisFPR=%xisCSR=%x use=%x\n    src2=ArchRegOperand: idx=%xrtype=%sisGPR=%xisFPR=%xisCSR=%x use=%x\n use=\n    imm=%x (usage=%s)\n  Control Flags:\n    ALU: AluCtrlFlags: isSub=%x isAdd=%x isSigned=%x logicOp=%s\n    Shift: ShiftCtrlFlags: isRight=%x isArithmetic=%x isRotate=%x isDoubleWord=%x\n    MulDiv: MulDivCtrlFlags: isDiv=%x isSigned=%x isWordOp=%x\n    Mem: MemCtrlFlags: size=%s isSignedLoad=%x isStore=%x isLoadLinked=%x isStoreCond=%x atomicOp=%x isFence=%x fenceMode=%x isCacheOp=%x cacheOpType=%x isPrefetch=%x\n    Branch: BranchCtrlFlags: condition=%s isJump=%x isLink=%x linkReg=ArchRegOperand: idx=%xrtype=%sisGPR=%xisFPR=%xisCSR=%x isIndirect=%x laCfIdx=%x\n    FPU: FpuCtrlFlags: opType=%x fpSizeSrc1=%s fpSizeSrc2=%s fpSizeDest=%s roundingMode=%x isIntegerDest=%x isSignedCvt=%x fmaNegSrc1=%x fcmpCond=%x\n    CSR: CsrCtrlFlags: csrAddr=%x isWrite=%x isRead=%x isExchange=%x useUimmAsSrc=%x\n    System: SystemCtrlFlags: sysCode=%x isExceptionReturn=%x isTlbOp=%x tlbOpType=%x\n  Status:\n    decodeEx=%s hasEx=%x\n    isMicrocode=%x entry=%x\n    isSerializing=%x isBranchOrJump=%x branchPrediction=BranchPredictionInfo: isTaken=%x target=%x wasPredicted=%x[0m", s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_pc, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isValid, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype_string, _zz_39, _zz_40, _zz_41, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype_string, _zz_42, _zz_43, _zz_44, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype_string, _zz_45, _zz_46, _zz_47, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_imm, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype_string, _zz_48, _zz_49, _zz_50, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode_string, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isSerializing, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target, s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted); // RenamePlugin.scala:L84
            end
          `endif
        `endif
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(((! s2_RobAlloc_isFiring) || RenamePlugin_logic_s2_logic_allocationOk)); // RenamePlugin.scala:L100
        `else
          if(!((! s2_RobAlloc_isFiring) || RenamePlugin_logic_s2_logic_allocationOk)) begin
            $display("FAILURE ASSERTION FAILED: Firing S2 stage with failed FreeList allocation!"); // RenamePlugin.scala:L100
            $finish;
          end
        `endif
      `endif
      if(FetchPipelinePlugin_doHardRedirect_listening) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LinkerPlugin.scala:L130
          `else
            if(!1'b0) begin
              $display("NOTE(LinkerPlugin.scala:130):  [normal] LinkerPlugin: Global doHardRedirect signal is asserted!"); // LinkerPlugin.scala:L130
            end
          `endif
        `endif
      end
      if(AluIntEU_AluIntEuPlugin_euInputPort_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LinkerPlugin.scala:L143
          `else
            if(!1'b0) begin
              $display("NOTE(LinkerPlugin.scala:143):  [normal] LinkerPlugin-Trace: Firing from IQ 'AluIntEU_IQ-0' to EU 'AluIntEU'. RobPtr=%x", AluIntEU_AluIntEuPlugin_euInputPort_payload_robPtr); // LinkerPlugin.scala:L143
            end
          `endif
        `endif
      end
      if(MulEU_MulEuPlugin_euInputPort_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LinkerPlugin.scala:L143
          `else
            if(!1'b0) begin
              $display("NOTE(LinkerPlugin.scala:143):  [normal] LinkerPlugin-Trace: Firing from IQ 'MulEU_IQ-1' to EU 'MulEU'. RobPtr=%x", MulEU_MulEuPlugin_euInputPort_payload_robPtr); // LinkerPlugin.scala:L143
            end
          `endif
        `endif
      end
      if(BranchEU_BranchEuPlugin_euInputPort_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LinkerPlugin.scala:L143
          `else
            if(!1'b0) begin
              $display("NOTE(LinkerPlugin.scala:143):  [normal] LinkerPlugin-Trace: Firing from IQ 'BranchEU_IQ-2' to EU 'BranchEU'. RobPtr=%x", BranchEU_BranchEuPlugin_euInputPort_payload_robPtr); // LinkerPlugin.scala:L143
            end
          `endif
        `endif
      end
      if(LsuEU_LsuEuPlugin_euInputPort_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LinkerPlugin.scala:L143
          `else
            if(!1'b0) begin
              $display("NOTE(LinkerPlugin.scala:143):  [normal] LinkerPlugin-Trace: Firing from IQ 'LsuEU_IQ-3' to EU 'LsuEU'. RobPtr=%x", LsuEU_LsuEuPlugin_euInputPort_payload_robPtr); // LinkerPlugin.scala:L143
            end
          `endif
        `endif
      end
      if(oneShot_20_io_pulseOut) begin
        if(when_Debug_l71_6) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_7};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_7); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(when_DispatchPlugin_l100) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // DispatchPlugin.scala:L101
          `else
            if(!1'b0) begin
              $display("NOTE(DispatchPlugin.scala:101):  [normal] DispatchPlugin: Firing robPtr=%x (UopCode=%s), s1_ready=%x, s2_ready=%x", s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr, s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode_string, DispatchPlugin_logic_src1InitialReady, DispatchPlugin_logic_src2InitialReady); // DispatchPlugin.scala:L101
            end
          `endif
        `endif
      end
      if(FetchPipelinePlugin_doHardRedirect_listening) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // DispatchPlugin.scala:L112
          `else
            if(!1'b0) begin
              $display("NOTE(DispatchPlugin.scala:112):  DispatchPlugin: (s3): Flushing pipeline due to hard redirect"); // DispatchPlugin.scala:L112
            end
          `endif
        `endif
      end
      if(DebugDisplayPlugin_logic_displayArea_divider_io_tick) begin
        DebugDisplayPlugin_logic_displayArea_dpToggle <= (! DebugDisplayPlugin_logic_displayArea_dpToggle);
      end
      if(s2_Execute_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // AluIntEuPlugin.scala:L107
          `else
            if(!1'b0) begin
              $display("NOTE(AluIntEuPlugin.scala:107):  [debug] [34mAluIntEu (AluIntEU) S2 Firing: RobPtr=%x, ResultData=%x, WritesPreg=%x, ImmUsage=%x, UseSrc2=%x op: AluCtrlFlags: isSub=%x isAdd=%x isSigned=%x logicOp=%s, lhs=%x, rhs=%x[0m", _zz_io_iqEntryIn_payload_robPtr, AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_data, AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_writesToPhysReg, _zz_51, _zz_io_iqEntryIn_payload_useSrc2, _zz_io_iqEntryIn_payload_aluCtrl_isSub, _zz_io_iqEntryIn_payload_aluCtrl_isAdd, _zz_io_iqEntryIn_payload_aluCtrl_isSigned, _zz_io_iqEntryIn_payload_aluCtrl_logicOp_string, _zz_io_iqEntryIn_payload_src1Data, _zz_io_iqEntryIn_payload_src2Data_1); // AluIntEuPlugin.scala:L107
            end
          `endif
        `endif
      end
      s1_ReadRegs_valid <= _zz_s1_ReadRegs_valid;
      if(when_Connection_l66_2) begin
        s1_ReadRegs_valid <= 1'b0;
      end
      s2_Execute_valid <= _zz_s2_Execute_valid;
      if(when_Connection_l66_1) begin
        s2_Execute_valid <= 1'b0;
      end
      s3_Writeback_valid <= _zz_s3_Writeback_valid;
      if(ROBPlugin_aggregatedFlushSignal_valid) begin
        s3_Writeback_valid <= 1'b0;
      end
      if(when_EuBasePlugin_l230) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L231
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:231):  EUBase (AluIntEU): Killing in-flight uop. robPtr=%x, flushTarget=%x", AluIntEU_AluIntEuPlugin_euResult_uop_robPtr, ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr); // EuBasePlugin.scala:L231
            end
          `endif
        `endif
      end
      if(AluIntEU_AluIntEuPlugin_euResult_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L243
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:243):  EUBase (AluIntEU): Result valid, writesToPreg=%x, hasException=%x, executionCompletes=%x, completesSuccessfully=%x, isFlushed=%x", AluIntEU_AluIntEuPlugin_euResult_writesToPreg, AluIntEU_AluIntEuPlugin_euResult_hasException, AluIntEU_AluIntEuPlugin_logicPhase_executionCompletes, AluIntEU_AluIntEuPlugin_logicPhase_completesSuccessfully, ROBPlugin_aggregatedFlushSignal_valid); // EuBasePlugin.scala:L243
            end
          `endif
        `endif
      end
      if(oneShot_21_io_pulseOut) begin
        if(when_Debug_l71_7) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_8};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_8); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(when_EuBasePlugin_l300) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L301
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:301):  [RAW_DEBUG] EU (AluIntEU) clearing BusyTable: physReg=%x, robPtr=%x", AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx, AluIntEU_AluIntEuPlugin_euResult_uop_robPtr); // EuBasePlugin.scala:L301
            end
          `endif
        `endif
      end
      if(mul_s2_Execute_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // MulEuPlugin.scala:L96
          `else
            if(!1'b0) begin
              $display("NOTE(MulEuPlugin.scala:96):  [normal] MulEuPlugin (MulEU) S2 Firing: RobPtr=%x, src1=%x, src2=%xmulDivCtrl=MulDivCtrlFlags: isDiv=%x isSigned=%x isWordOp=%x", _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_6, _zz_A, _zz_B, _zz_23, _zz_24, _zz_25); // MulEuPlugin.scala:L96
            end
          `endif
        `endif
      end
      if(mul_s7_Writeback_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // MulEuPlugin.scala:L114
          `else
            if(!1'b0) begin
              $display("NOTE(MulEuPlugin.scala:114):  [normal] MulEuPlugin (MulEU) S7 Firing: RobPtr=%x, Result=%xmulDivCtrl=MulDivCtrlFlags: isDiv=%x isSigned=%x isWordOp=%x", _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_5, _zz_MulEU_MulEuPlugin_euResult_data, _zz_20, _zz_21, _zz_22); // MulEuPlugin.scala:L114
            end
          `endif
        `endif
      end
      mul_s1_ReadRegs_valid <= _zz_mul_s1_ReadRegs_valid;
      if(when_Connection_l66_8) begin
        mul_s1_ReadRegs_valid <= 1'b0;
      end
      mul_s2_Execute_valid <= _zz_mul_s2_Execute_valid;
      if(when_Connection_l66_7) begin
        mul_s2_Execute_valid <= 1'b0;
      end
      mul_s3_Execute_valid <= _zz_mul_s3_Execute_valid;
      if(when_Connection_l66_6) begin
        mul_s3_Execute_valid <= 1'b0;
      end
      mul_s4_Execute_valid <= _zz_mul_s4_Execute_valid;
      if(when_Connection_l66_5) begin
        mul_s4_Execute_valid <= 1'b0;
      end
      mul_s5_Execute_valid <= _zz_mul_s5_Execute_valid;
      if(when_Connection_l66_4) begin
        mul_s5_Execute_valid <= 1'b0;
      end
      mul_s6_Execute_valid <= _zz_mul_s6_Execute_valid;
      if(when_Connection_l66_3) begin
        mul_s6_Execute_valid <= 1'b0;
      end
      mul_s7_Writeback_valid <= _zz_mul_s7_Writeback_valid;
      if(ROBPlugin_aggregatedFlushSignal_valid) begin
        mul_s7_Writeback_valid <= 1'b0;
      end
      if(when_EuBasePlugin_l230_1) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L231
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:231):  EUBase (MulEU): Killing in-flight uop. robPtr=%x, flushTarget=%x", MulEU_MulEuPlugin_euResult_uop_robPtr, ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr); // EuBasePlugin.scala:L231
            end
          `endif
        `endif
      end
      if(MulEU_MulEuPlugin_euResult_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L243
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:243):  EUBase (MulEU): Result valid, writesToPreg=%x, hasException=%x, executionCompletes=%x, completesSuccessfully=%x, isFlushed=%x", MulEU_MulEuPlugin_euResult_writesToPreg, MulEU_MulEuPlugin_euResult_hasException, MulEU_MulEuPlugin_logicPhase_executionCompletes, MulEU_MulEuPlugin_logicPhase_completesSuccessfully, ROBPlugin_aggregatedFlushSignal_valid); // EuBasePlugin.scala:L243
            end
          `endif
        `endif
      end
      if(oneShot_22_io_pulseOut) begin
        if(when_Debug_l71_8) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_9};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_9); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(when_EuBasePlugin_l300_1) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L301
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:301):  [RAW_DEBUG] EU (MulEU) clearing BusyTable: physReg=%x, robPtr=%x", MulEU_MulEuPlugin_euResult_uop_physDest_idx, MulEU_MulEuPlugin_euResult_uop_robPtr); // EuBasePlugin.scala:L301
            end
          `endif
        `endif
      end
      if(s0_Dispatch_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BranchEuPlugin.scala:L98
          `else
            if(!1'b0) begin
              $display("NOTE(BranchEuPlugin.scala:98):  [BranchEU-S0] DISPATCH: PC=0x%x", _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_3); // BranchEuPlugin.scala:L98
            end
          `endif
        `endif
      end
      if(s1_Calc_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BranchEuPlugin.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(BranchEuPlugin.scala:104):  [BranchEU-S1-Calc] CALC START: PC=0x%x", _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_2); // BranchEuPlugin.scala:L104
            end
          `endif
        `endif
      end
      if(s2_Select_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BranchEuPlugin.scala:L151
          `else
            if(!1'b0) begin
              $display("NOTE(BranchEuPlugin.scala:151):  [BranchEU-S2-Select] SELECT START: PC=0x%x, branchTaken(from S1)=%x", _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_1, _zz_BranchEU_BranchEuPlugin_euResult_data_2); // BranchEuPlugin.scala:L151
            end
          `endif
        `endif
      end
      if(s2_Select_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BranchEuPlugin.scala:L191
          `else
            if(!1'b0) begin
              $display("NOTE(BranchEuPlugin.scala:191):  [BranchEU-S2-Select] PREDICTION: wasPredicted(valid)=%x: predictedTaken=%x, actuallyTaken=%x, finalTarget=0x%x, mispredicted=%x", _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted_1, _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken_1, _zz_BranchEU_BranchEuPlugin_euResult_isTaken_1, _zz_BranchEU_BranchEuPlugin_euResult_data_6, _zz_52); // BranchEuPlugin.scala:L191
            end
          `endif
        `endif
      end
      if(s3_Result_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BranchEuPlugin.scala:L226
          `else
            if(!1'b0) begin
              $display("NOTE(BranchEuPlugin.scala:226):  [BranchEU-S3-Result] RESULT: euResult.valid=1, writesToPreg=%x, data=0x%x, mispredicted=%x", BranchEU_BranchEuPlugin_euResult_writesToPreg, BranchEU_BranchEuPlugin_euResult_data, BranchEU_BranchEuPlugin_euResult_isMispredictedBranch); // BranchEuPlugin.scala:L226
            end
          `endif
        `endif
      end
      s1_Calc_valid <= _zz_s1_Calc_valid;
      if(when_Connection_l66_10) begin
        s1_Calc_valid <= 1'b0;
      end
      s2_Select_valid <= _zz_s2_Select_valid;
      if(when_Connection_l66_9) begin
        s2_Select_valid <= 1'b0;
      end
      s3_Result_valid <= _zz_s3_Result_valid;
      if(ROBPlugin_aggregatedFlushSignal_valid) begin
        s3_Result_valid <= 1'b0;
      end
      if(when_EuBasePlugin_l230_2) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L231
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:231):  EUBase (BranchEU): Killing in-flight uop. robPtr=%x, flushTarget=%x", BranchEU_BranchEuPlugin_euResult_uop_robPtr, ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr); // EuBasePlugin.scala:L231
            end
          `endif
        `endif
      end
      if(BranchEU_BranchEuPlugin_euResult_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L243
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:243):  EUBase (BranchEU): Result valid, writesToPreg=%x, hasException=%x, executionCompletes=%x, completesSuccessfully=%x, isFlushed=%x", BranchEU_BranchEuPlugin_euResult_writesToPreg, BranchEU_BranchEuPlugin_euResult_hasException, BranchEU_BranchEuPlugin_logicPhase_executionCompletes, BranchEU_BranchEuPlugin_logicPhase_completesSuccessfully, ROBPlugin_aggregatedFlushSignal_valid); // EuBasePlugin.scala:L243
            end
          `endif
        `endif
      end
      if(oneShot_23_io_pulseOut) begin
        if(when_Debug_l71_9) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_10};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_10); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(when_EuBasePlugin_l300_2) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L301
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:301):  [RAW_DEBUG] EU (BranchEU) clearing BusyTable: physReg=%x, robPtr=%x", BranchEU_BranchEuPlugin_euResult_uop_physDest_idx, BranchEU_BranchEuPlugin_euResult_uop_robPtr); // EuBasePlugin.scala:L301
            end
          `endif
        `endif
      end
      if(when_LsuEuPlugin_l141) begin
        if(LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // LsuEuPlugin.scala:L142
            `else
              if(!1'b0) begin
                $display("NOTE(LsuEuPlugin.scala:142):  [normal] [LsuEu] Dispatched LOAD to LQ: robPtr=%x", LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr); // LsuEuPlugin.scala:L142
              end
            `endif
          `endif
        end
        if(LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isStore) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // LsuEuPlugin.scala:L143
            `else
              if(!1'b0) begin
                $display("NOTE(LsuEuPlugin.scala:143):  [normal] [LsuEu] Dispatched STORE to SB: robPtr=%x", LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr); // LsuEuPlugin.scala:L143
              end
            `endif
          `endif
        end
      end
      if(when_EuBasePlugin_l230_3) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L231
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:231):  EUBase (LsuEU): Killing in-flight uop. robPtr=%x, flushTarget=%x", LsuEU_LsuEuPlugin_euResult_uop_robPtr, ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr); // EuBasePlugin.scala:L231
            end
          `endif
        `endif
      end
      if(LsuEU_LsuEuPlugin_euResult_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L243
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:243):  EUBase (LsuEU): Result valid, writesToPreg=%x, hasException=%x, executionCompletes=%x, completesSuccessfully=%x, isFlushed=%x", LsuEU_LsuEuPlugin_euResult_writesToPreg, LsuEU_LsuEuPlugin_euResult_hasException, LsuEU_LsuEuPlugin_logicPhase_executionCompletes, LsuEU_LsuEuPlugin_logicPhase_completesSuccessfully, ROBPlugin_aggregatedFlushSignal_valid); // EuBasePlugin.scala:L243
            end
          `endif
        `endif
      end
      if(oneShot_24_io_pulseOut) begin
        if(when_Debug_l71_10) begin
          _zz_when_Debug_l71 <= {3'd0, _zz_when_Debug_l71_11};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_11); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(when_EuBasePlugin_l300_3) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // EuBasePlugin.scala:L301
          `else
            if(!1'b0) begin
              $display("NOTE(EuBasePlugin.scala:301):  [RAW_DEBUG] EU (LsuEU) clearing BusyTable: physReg=%x, robPtr=%x", LsuEU_LsuEuPlugin_euResult_uop_physDest_idx, LsuEU_LsuEuPlugin_euResult_uop_robPtr); // EuBasePlugin.scala:L301
            end
          `endif
        `endif
      end
      if(s0_Decode_ready_output) begin
        s1_Rename_valid <= _zz_s1_Rename_valid;
      end
      if(when_Connection_l66_11) begin
        s1_Rename_valid <= 1'b0;
      end
      if(s1_Rename_ready_output) begin
        s2_RobAlloc_valid <= _zz_s2_RobAlloc_valid;
      end
      if(when_Connection_l66) begin
        s2_RobAlloc_valid <= 1'b0;
      end
      if(s2_RobAlloc_ready_output) begin
        s3_Dispatch_valid <= _zz_s3_Dispatch_valid;
      end
      if(when_Connection_l66) begin
        s3_Dispatch_valid <= 1'b0;
      end
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid;
      if(LsuEU_LsuEuPlugin_hw_aguPort_flush) begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid <= 1'b0;
      end
      if(_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // AddressGenerationUnit.scala:L266
          `else
            if(!1'b0) begin
              $display("NOTE(AddressGenerationUnit.scala:266):  [normal] [AGU-0-S1-Output-Debug] s1.payload=AguInput(qPtr=%x,basePhysReg=%x,immediate=%x,accessSize=%s,usePc=%x,pc=%x,dataReg=%x,robPtr=%x,isLoad=%x,isStore=%x,isFlush=%x,isIO=%x,physDst=%x) baseData=0x%x ==> effAddr=0x%x", _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr, _zz_when_AddressGenerationUnit_l215, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_string, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc, _zz_when_AddressGenerationUnit_l220, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad, _zz_when_AddressGenerationUnit_l220_1, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_3, _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_4); // AddressGenerationUnit.scala:L266
            end
          `endif
        `endif
      end
      if(_zz_LsuEU_LsuEuPlugin_hw_aguPort_input_ready) begin
        _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid_2 <= (_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_valid && (! LsuEU_LsuEuPlugin_hw_aguPort_flush));
      end
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_valid <= LoadQueuePlugin_logic_loadQueue_completionInfo_valid;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromFwd <= LoadQueuePlugin_logic_loadQueue_completionInfo_fromFwd;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromDCache <= LoadQueuePlugin_logic_loadQueue_completionInfo_fromDCache;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromMMIO <= LoadQueuePlugin_logic_loadQueue_completionInfo_fromMMIO;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_fromEarlyExc <= LoadQueuePlugin_logic_loadQueue_completionInfo_fromEarlyExc;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_data <= LoadQueuePlugin_logic_loadQueue_completionInfo_data;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_hasFault <= LoadQueuePlugin_logic_loadQueue_completionInfo_hasFault;
      LoadQueuePlugin_logic_loadQueue_completionInfoReg_exceptionCode <= LoadQueuePlugin_logic_loadQueue_completionInfo_exceptionCode;
      LoadQueuePlugin_logic_loadQueue_sbQueryRspValid <= StoreBufferPlugin_hw_sqQueryPort_cmd_valid;
      LoadQueuePlugin_logic_loadQueue_registeredFlush_valid <= LoadQueuePlugin_logic_loadQueue_flushInProgress;
      LoadQueuePlugin_logic_loadQueue_registeredFlush_targetRobPtr <= ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr;
      if(LoadQueuePlugin_logic_pushCmd_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L304
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:304):  [normal] [LQ] PUSH from LsuEu: robPtr=%x addr=%x to slotIdx=%x", LoadQueuePlugin_logic_pushCmd_payload_robPtr, LoadQueuePlugin_logic_pushCmd_payload_address, LoadQueuePlugin_logic_loadQueue_pushIdx); // LoadQueuePlugin.scala:L304
            end
          `endif
        `endif
      end
      if(StoreBufferPlugin_hw_sqQueryPort_cmd_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L326
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:326):  [normal] [LQ-Fwd] QUERY: robPtr=%x addr=%x", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr, LoadQueuePlugin_logic_loadQueue_slots_0_address); // LoadQueuePlugin.scala:L326
            end
          `endif
        `endif
      end
      if(when_LoadQueuePlugin_l329) begin
        if(LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_hit) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // LoadQueuePlugin.scala:L334
            `else
              if(!1'b0) begin
                $display("NOTE(LoadQueuePlugin.scala:334):  [normal] [LQ-Fwd] HIT: robPtr=%x, data=%x. Will complete via popOnFwdHit.", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr, LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_data); // LoadQueuePlugin.scala:L334
              end
            `endif
          `endif
        end else begin
          if(when_LoadQueuePlugin_l335) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // LoadQueuePlugin.scala:L336
              `else
                if(!1'b0) begin
                  $display("NOTE(LoadQueuePlugin.scala:336):  [normal] [LQ-Fwd] STALL: robPtr=%x has dependency...", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr); // LoadQueuePlugin.scala:L336
                end
              `endif
            `endif
          end else begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // LoadQueuePlugin.scala:L339
              `else
                if(!1'b0) begin
                  $display("NOTE(LoadQueuePlugin.scala:339):  [normal] [LQ-Fwd] MISS: robPtr=%x is clear to access D-Cache or MMIO.", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr); // LoadQueuePlugin.scala:L339
                end
              `endif
            `endif
          end
        end
      end
      if(when_LoadQueuePlugin_l350) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L352
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:352):  [normal] [LQ] Early exception for robPtr=%x, marking ready for exception handling", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr); // LoadQueuePlugin.scala:L352
            end
          `endif
        `endif
      end
      if(LoadQueuePlugin_hw_dCacheLoadPort_cmd_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L377
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:377):  [normal] [LQ-DCache] SEND_TO_DCACHE: robPtr=%x addr=%x", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr, LoadQueuePlugin_logic_loadQueue_slots_0_address); // LoadQueuePlugin.scala:L377
            end
          `endif
        `endif
      end
      if(LoadQueuePlugin_logic_loadQueue_mmioCmdFired) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L392
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:392):  [normal] [LQ-MMIO] SEND_TO_MMIO: robPtr=%x addr=%x", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr, LoadQueuePlugin_logic_loadQueue_slots_0_address); // LoadQueuePlugin.scala:L392
            end
          `endif
        `endif
      end
      if(when_LoadQueuePlugin_l409) begin
        if(LoadQueuePlugin_hw_dCacheLoadPort_rsp_payload_redo) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // LoadQueuePlugin.scala:L413
            `else
              if(!1'b0) begin
                $display("NOTE(LoadQueuePlugin.scala:413):  [normal] [LQ-DCache] REDO received for robPtr=%x", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr); // LoadQueuePlugin.scala:L413
              end
            `endif
          `endif
        end
      end
      if(when_LoadQueuePlugin_l508) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L511
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:511):  [normal] [LQ] FLUSH (Exec): Invalidating slotIdx=0 (robPtr=%x)", LoadQueuePlugin_logic_loadQueue_slots_0_robPtr); // LoadQueuePlugin.scala:L511
            end
          `endif
        `endif
      end
      if(when_LoadQueuePlugin_l508_1) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L511
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:511):  [normal] [LQ] FLUSH (Exec): Invalidating slotIdx=1 (robPtr=%x)", LoadQueuePlugin_logic_loadQueue_slots_1_robPtr); // LoadQueuePlugin.scala:L511
            end
          `endif
        `endif
      end
      if(when_LoadQueuePlugin_l508_2) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L511
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:511):  [normal] [LQ] FLUSH (Exec): Invalidating slotIdx=2 (robPtr=%x)", LoadQueuePlugin_logic_loadQueue_slots_2_robPtr); // LoadQueuePlugin.scala:L511
            end
          `endif
        `endif
      end
      if(when_LoadQueuePlugin_l508_3) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // LoadQueuePlugin.scala:L511
          `else
            if(!1'b0) begin
              $display("NOTE(LoadQueuePlugin.scala:511):  [normal] [LQ] FLUSH (Exec): Invalidating slotIdx=3 (robPtr=%x)", LoadQueuePlugin_logic_loadQueue_slots_3_robPtr); // LoadQueuePlugin.scala:L511
            end
          `endif
        `endif
      end
      LoadQueuePlugin_logic_loadQueue_slots_0_valid <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_valid;
      LoadQueuePlugin_logic_loadQueue_slots_0_address <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_address;
      LoadQueuePlugin_logic_loadQueue_slots_0_size <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_size;
      LoadQueuePlugin_logic_loadQueue_slots_0_robPtr <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_robPtr;
      LoadQueuePlugin_logic_loadQueue_slots_0_pdest <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_pdest;
      LoadQueuePlugin_logic_loadQueue_slots_0_isIO <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_isIO;
      LoadQueuePlugin_logic_loadQueue_slots_0_hasException <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_hasException;
      LoadQueuePlugin_logic_loadQueue_slots_0_exceptionCode <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_exceptionCode;
      LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForFwdRsp;
      LoadQueuePlugin_logic_loadQueue_slots_0_isStalledByDependency <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_isStalledByDependency;
      LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_isReadyForDCache;
      LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp <= LoadQueuePlugin_logic_loadQueue_slotsNext_0_isWaitingForRsp;
      LoadQueuePlugin_logic_loadQueue_slots_1_valid <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_valid;
      LoadQueuePlugin_logic_loadQueue_slots_1_address <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_address;
      LoadQueuePlugin_logic_loadQueue_slots_1_size <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_size;
      LoadQueuePlugin_logic_loadQueue_slots_1_robPtr <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_robPtr;
      LoadQueuePlugin_logic_loadQueue_slots_1_pdest <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_pdest;
      LoadQueuePlugin_logic_loadQueue_slots_1_isIO <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_isIO;
      LoadQueuePlugin_logic_loadQueue_slots_1_hasException <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_hasException;
      LoadQueuePlugin_logic_loadQueue_slots_1_exceptionCode <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_exceptionCode;
      LoadQueuePlugin_logic_loadQueue_slots_1_isWaitingForFwdRsp <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForFwdRsp;
      LoadQueuePlugin_logic_loadQueue_slots_1_isStalledByDependency <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_isStalledByDependency;
      LoadQueuePlugin_logic_loadQueue_slots_1_isReadyForDCache <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_isReadyForDCache;
      LoadQueuePlugin_logic_loadQueue_slots_1_isWaitingForRsp <= LoadQueuePlugin_logic_loadQueue_slotsNext_1_isWaitingForRsp;
      LoadQueuePlugin_logic_loadQueue_slots_2_valid <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_valid;
      LoadQueuePlugin_logic_loadQueue_slots_2_address <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_address;
      LoadQueuePlugin_logic_loadQueue_slots_2_size <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_size;
      LoadQueuePlugin_logic_loadQueue_slots_2_robPtr <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_robPtr;
      LoadQueuePlugin_logic_loadQueue_slots_2_pdest <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_pdest;
      LoadQueuePlugin_logic_loadQueue_slots_2_isIO <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_isIO;
      LoadQueuePlugin_logic_loadQueue_slots_2_hasException <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_hasException;
      LoadQueuePlugin_logic_loadQueue_slots_2_exceptionCode <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_exceptionCode;
      LoadQueuePlugin_logic_loadQueue_slots_2_isWaitingForFwdRsp <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForFwdRsp;
      LoadQueuePlugin_logic_loadQueue_slots_2_isStalledByDependency <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_isStalledByDependency;
      LoadQueuePlugin_logic_loadQueue_slots_2_isReadyForDCache <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_isReadyForDCache;
      LoadQueuePlugin_logic_loadQueue_slots_2_isWaitingForRsp <= LoadQueuePlugin_logic_loadQueue_slotsNext_2_isWaitingForRsp;
      LoadQueuePlugin_logic_loadQueue_slots_3_valid <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_valid;
      LoadQueuePlugin_logic_loadQueue_slots_3_address <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_address;
      LoadQueuePlugin_logic_loadQueue_slots_3_size <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_size;
      LoadQueuePlugin_logic_loadQueue_slots_3_robPtr <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_robPtr;
      LoadQueuePlugin_logic_loadQueue_slots_3_pdest <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_pdest;
      LoadQueuePlugin_logic_loadQueue_slots_3_isIO <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_isIO;
      LoadQueuePlugin_logic_loadQueue_slots_3_hasException <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_hasException;
      LoadQueuePlugin_logic_loadQueue_slots_3_exceptionCode <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_exceptionCode;
      LoadQueuePlugin_logic_loadQueue_slots_3_isWaitingForFwdRsp <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForFwdRsp;
      LoadQueuePlugin_logic_loadQueue_slots_3_isStalledByDependency <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_isStalledByDependency;
      LoadQueuePlugin_logic_loadQueue_slots_3_isReadyForDCache <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_isReadyForDCache;
      LoadQueuePlugin_logic_loadQueue_slots_3_isWaitingForRsp <= LoadQueuePlugin_logic_loadQueue_slotsNext_3_isWaitingForRsp;
      if(AluIntEU_AluIntEuPlugin_gprReadPorts_0_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:104):  [normal] [PRegPlugin] Read from reg[%x] -> %x", AluIntEU_AluIntEuPlugin_gprReadPorts_0_address, AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp); // PhysicalRegFile.scala:L104
            end
          `endif
        `endif
      end
      if(AluIntEU_AluIntEuPlugin_gprReadPorts_1_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:104):  [normal] [PRegPlugin] Read from reg[%x] -> %x", AluIntEU_AluIntEuPlugin_gprReadPorts_1_address, AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp); // PhysicalRegFile.scala:L104
            end
          `endif
        `endif
      end
      if(MulEU_MulEuPlugin_gprReadPorts_0_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:104):  [normal] [PRegPlugin] Read from reg[%x] -> %x", MulEU_MulEuPlugin_gprReadPorts_0_address, MulEU_MulEuPlugin_gprReadPorts_0_rsp); // PhysicalRegFile.scala:L104
            end
          `endif
        `endif
      end
      if(MulEU_MulEuPlugin_gprReadPorts_1_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:104):  [normal] [PRegPlugin] Read from reg[%x] -> %x", MulEU_MulEuPlugin_gprReadPorts_1_address, MulEU_MulEuPlugin_gprReadPorts_1_rsp); // PhysicalRegFile.scala:L104
            end
          `endif
        `endif
      end
      if(BranchEU_BranchEuPlugin_gprReadPorts_0_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:104):  [normal] [PRegPlugin] Read from reg[%x] -> %x", BranchEU_BranchEuPlugin_gprReadPorts_0_address, BranchEU_BranchEuPlugin_gprReadPorts_0_rsp); // PhysicalRegFile.scala:L104
            end
          `endif
        `endif
      end
      if(BranchEU_BranchEuPlugin_gprReadPorts_1_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:104):  [normal] [PRegPlugin] Read from reg[%x] -> %x", BranchEU_BranchEuPlugin_gprReadPorts_1_address, BranchEU_BranchEuPlugin_gprReadPorts_1_rsp); // PhysicalRegFile.scala:L104
            end
          `endif
        `endif
      end
      if(LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:104):  [normal] [PRegPlugin] Read from reg[%x] -> %x", LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_address, LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp); // PhysicalRegFile.scala:L104
            end
          `endif
        `endif
      end
      if(LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L104
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:104):  [normal] [PRegPlugin] Read from reg[%x] -> %x", LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_address, LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp); // PhysicalRegFile.scala:L104
            end
          `endif
        `endif
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((AluIntEU_AluIntEuPlugin_gprWritePort_valid && MulEU_MulEuPlugin_gprWritePort_valid) && (AluIntEU_AluIntEuPlugin_gprWritePort_address == MulEU_MulEuPlugin_gprWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((AluIntEU_AluIntEuPlugin_gprWritePort_valid && MulEU_MulEuPlugin_gprWritePort_valid) && (AluIntEU_AluIntEuPlugin_gprWritePort_address == MulEU_MulEuPlugin_gprWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between AluIntEU.gprWritePort and MulEU.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((AluIntEU_AluIntEuPlugin_gprWritePort_valid && BranchEU_BranchEuPlugin_gprWritePort_valid) && (AluIntEU_AluIntEuPlugin_gprWritePort_address == BranchEU_BranchEuPlugin_gprWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((AluIntEU_AluIntEuPlugin_gprWritePort_valid && BranchEU_BranchEuPlugin_gprWritePort_valid) && (AluIntEU_AluIntEuPlugin_gprWritePort_address == BranchEU_BranchEuPlugin_gprWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between AluIntEU.gprWritePort and BranchEU.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((AluIntEU_AluIntEuPlugin_gprWritePort_valid && LsuEU_LsuEuPlugin_gprWritePort_valid) && (AluIntEU_AluIntEuPlugin_gprWritePort_address == LsuEU_LsuEuPlugin_gprWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((AluIntEU_AluIntEuPlugin_gprWritePort_valid && LsuEU_LsuEuPlugin_gprWritePort_valid) && (AluIntEU_AluIntEuPlugin_gprWritePort_address == LsuEU_LsuEuPlugin_gprWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between AluIntEU.gprWritePort and LsuEU.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((AluIntEU_AluIntEuPlugin_gprWritePort_valid && LoadQueuePlugin_hw_prfWritePort_valid) && (AluIntEU_AluIntEuPlugin_gprWritePort_address == LoadQueuePlugin_hw_prfWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((AluIntEU_AluIntEuPlugin_gprWritePort_valid && LoadQueuePlugin_hw_prfWritePort_valid) && (AluIntEU_AluIntEuPlugin_gprWritePort_address == LoadQueuePlugin_hw_prfWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between AluIntEU.gprWritePort and LQ.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((MulEU_MulEuPlugin_gprWritePort_valid && BranchEU_BranchEuPlugin_gprWritePort_valid) && (MulEU_MulEuPlugin_gprWritePort_address == BranchEU_BranchEuPlugin_gprWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((MulEU_MulEuPlugin_gprWritePort_valid && BranchEU_BranchEuPlugin_gprWritePort_valid) && (MulEU_MulEuPlugin_gprWritePort_address == BranchEU_BranchEuPlugin_gprWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between MulEU.gprWritePort and BranchEU.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((MulEU_MulEuPlugin_gprWritePort_valid && LsuEU_LsuEuPlugin_gprWritePort_valid) && (MulEU_MulEuPlugin_gprWritePort_address == LsuEU_LsuEuPlugin_gprWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((MulEU_MulEuPlugin_gprWritePort_valid && LsuEU_LsuEuPlugin_gprWritePort_valid) && (MulEU_MulEuPlugin_gprWritePort_address == LsuEU_LsuEuPlugin_gprWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between MulEU.gprWritePort and LsuEU.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((MulEU_MulEuPlugin_gprWritePort_valid && LoadQueuePlugin_hw_prfWritePort_valid) && (MulEU_MulEuPlugin_gprWritePort_address == LoadQueuePlugin_hw_prfWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((MulEU_MulEuPlugin_gprWritePort_valid && LoadQueuePlugin_hw_prfWritePort_valid) && (MulEU_MulEuPlugin_gprWritePort_address == LoadQueuePlugin_hw_prfWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between MulEU.gprWritePort and LQ.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((BranchEU_BranchEuPlugin_gprWritePort_valid && LsuEU_LsuEuPlugin_gprWritePort_valid) && (BranchEU_BranchEuPlugin_gprWritePort_address == LsuEU_LsuEuPlugin_gprWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((BranchEU_BranchEuPlugin_gprWritePort_valid && LsuEU_LsuEuPlugin_gprWritePort_valid) && (BranchEU_BranchEuPlugin_gprWritePort_address == LsuEU_LsuEuPlugin_gprWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between BranchEU.gprWritePort and LsuEU.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((BranchEU_BranchEuPlugin_gprWritePort_valid && LoadQueuePlugin_hw_prfWritePort_valid) && (BranchEU_BranchEuPlugin_gprWritePort_address == LoadQueuePlugin_hw_prfWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((BranchEU_BranchEuPlugin_gprWritePort_valid && LoadQueuePlugin_hw_prfWritePort_valid) && (BranchEU_BranchEuPlugin_gprWritePort_address == LoadQueuePlugin_hw_prfWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between BranchEU.gprWritePort and LQ.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((LsuEU_LsuEuPlugin_gprWritePort_valid && LoadQueuePlugin_hw_prfWritePort_valid) && (LsuEU_LsuEuPlugin_gprWritePort_address == LoadQueuePlugin_hw_prfWritePort_address)))); // PhysicalRegFile.scala:L118
        `else
          if(!(! ((LsuEU_LsuEuPlugin_gprWritePort_valid && LoadQueuePlugin_hw_prfWritePort_valid) && (LsuEU_LsuEuPlugin_gprWritePort_address == LoadQueuePlugin_hw_prfWritePort_address)))) begin
            $display("FAILURE CRITICAL ERROR: Concurrent write to the same physical register detected between LsuEU.gprWritePort and LQ.gprWritePort. This is a design flaw in the pipeline scheduling logic."); // PhysicalRegFile.scala:L118
            $finish;
          end
        `endif
      `endif
      if(when_PhysicalRegFile_l130) begin
        if(_zz_58[0]) begin
          PhysicalRegFilePlugin_logic_regFile_0 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[1]) begin
          PhysicalRegFilePlugin_logic_regFile_1 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[2]) begin
          PhysicalRegFilePlugin_logic_regFile_2 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[3]) begin
          PhysicalRegFilePlugin_logic_regFile_3 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[4]) begin
          PhysicalRegFilePlugin_logic_regFile_4 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[5]) begin
          PhysicalRegFilePlugin_logic_regFile_5 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[6]) begin
          PhysicalRegFilePlugin_logic_regFile_6 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[7]) begin
          PhysicalRegFilePlugin_logic_regFile_7 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[8]) begin
          PhysicalRegFilePlugin_logic_regFile_8 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[9]) begin
          PhysicalRegFilePlugin_logic_regFile_9 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[10]) begin
          PhysicalRegFilePlugin_logic_regFile_10 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[11]) begin
          PhysicalRegFilePlugin_logic_regFile_11 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[12]) begin
          PhysicalRegFilePlugin_logic_regFile_12 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[13]) begin
          PhysicalRegFilePlugin_logic_regFile_13 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[14]) begin
          PhysicalRegFilePlugin_logic_regFile_14 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[15]) begin
          PhysicalRegFilePlugin_logic_regFile_15 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[16]) begin
          PhysicalRegFilePlugin_logic_regFile_16 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[17]) begin
          PhysicalRegFilePlugin_logic_regFile_17 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[18]) begin
          PhysicalRegFilePlugin_logic_regFile_18 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[19]) begin
          PhysicalRegFilePlugin_logic_regFile_19 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[20]) begin
          PhysicalRegFilePlugin_logic_regFile_20 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[21]) begin
          PhysicalRegFilePlugin_logic_regFile_21 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[22]) begin
          PhysicalRegFilePlugin_logic_regFile_22 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[23]) begin
          PhysicalRegFilePlugin_logic_regFile_23 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[24]) begin
          PhysicalRegFilePlugin_logic_regFile_24 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[25]) begin
          PhysicalRegFilePlugin_logic_regFile_25 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[26]) begin
          PhysicalRegFilePlugin_logic_regFile_26 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[27]) begin
          PhysicalRegFilePlugin_logic_regFile_27 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[28]) begin
          PhysicalRegFilePlugin_logic_regFile_28 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[29]) begin
          PhysicalRegFilePlugin_logic_regFile_29 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[30]) begin
          PhysicalRegFilePlugin_logic_regFile_30 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[31]) begin
          PhysicalRegFilePlugin_logic_regFile_31 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[32]) begin
          PhysicalRegFilePlugin_logic_regFile_32 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[33]) begin
          PhysicalRegFilePlugin_logic_regFile_33 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[34]) begin
          PhysicalRegFilePlugin_logic_regFile_34 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[35]) begin
          PhysicalRegFilePlugin_logic_regFile_35 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[36]) begin
          PhysicalRegFilePlugin_logic_regFile_36 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[37]) begin
          PhysicalRegFilePlugin_logic_regFile_37 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[38]) begin
          PhysicalRegFilePlugin_logic_regFile_38 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[39]) begin
          PhysicalRegFilePlugin_logic_regFile_39 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[40]) begin
          PhysicalRegFilePlugin_logic_regFile_40 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[41]) begin
          PhysicalRegFilePlugin_logic_regFile_41 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[42]) begin
          PhysicalRegFilePlugin_logic_regFile_42 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[43]) begin
          PhysicalRegFilePlugin_logic_regFile_43 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[44]) begin
          PhysicalRegFilePlugin_logic_regFile_44 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[45]) begin
          PhysicalRegFilePlugin_logic_regFile_45 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[46]) begin
          PhysicalRegFilePlugin_logic_regFile_46 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[47]) begin
          PhysicalRegFilePlugin_logic_regFile_47 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[48]) begin
          PhysicalRegFilePlugin_logic_regFile_48 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[49]) begin
          PhysicalRegFilePlugin_logic_regFile_49 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[50]) begin
          PhysicalRegFilePlugin_logic_regFile_50 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[51]) begin
          PhysicalRegFilePlugin_logic_regFile_51 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[52]) begin
          PhysicalRegFilePlugin_logic_regFile_52 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[53]) begin
          PhysicalRegFilePlugin_logic_regFile_53 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[54]) begin
          PhysicalRegFilePlugin_logic_regFile_54 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[55]) begin
          PhysicalRegFilePlugin_logic_regFile_55 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[56]) begin
          PhysicalRegFilePlugin_logic_regFile_56 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[57]) begin
          PhysicalRegFilePlugin_logic_regFile_57 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[58]) begin
          PhysicalRegFilePlugin_logic_regFile_58 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[59]) begin
          PhysicalRegFilePlugin_logic_regFile_59 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[60]) begin
          PhysicalRegFilePlugin_logic_regFile_60 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[61]) begin
          PhysicalRegFilePlugin_logic_regFile_61 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[62]) begin
          PhysicalRegFilePlugin_logic_regFile_62 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        if(_zz_58[63]) begin
          PhysicalRegFilePlugin_logic_regFile_63 <= AluIntEU_AluIntEuPlugin_gprWritePort_data;
        end
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L134
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:134):  [normal] [PRegPlugin] Write from `AluIntEU.gprWritePort` to reg[%x] with data %x", AluIntEU_AluIntEuPlugin_gprWritePort_address, AluIntEU_AluIntEuPlugin_gprWritePort_data); // PhysicalRegFile.scala:L134
            end
          `endif
        `endif
      end
      if(when_PhysicalRegFile_l130_1) begin
        if(_zz_59[0]) begin
          PhysicalRegFilePlugin_logic_regFile_0 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[1]) begin
          PhysicalRegFilePlugin_logic_regFile_1 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[2]) begin
          PhysicalRegFilePlugin_logic_regFile_2 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[3]) begin
          PhysicalRegFilePlugin_logic_regFile_3 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[4]) begin
          PhysicalRegFilePlugin_logic_regFile_4 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[5]) begin
          PhysicalRegFilePlugin_logic_regFile_5 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[6]) begin
          PhysicalRegFilePlugin_logic_regFile_6 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[7]) begin
          PhysicalRegFilePlugin_logic_regFile_7 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[8]) begin
          PhysicalRegFilePlugin_logic_regFile_8 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[9]) begin
          PhysicalRegFilePlugin_logic_regFile_9 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[10]) begin
          PhysicalRegFilePlugin_logic_regFile_10 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[11]) begin
          PhysicalRegFilePlugin_logic_regFile_11 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[12]) begin
          PhysicalRegFilePlugin_logic_regFile_12 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[13]) begin
          PhysicalRegFilePlugin_logic_regFile_13 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[14]) begin
          PhysicalRegFilePlugin_logic_regFile_14 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[15]) begin
          PhysicalRegFilePlugin_logic_regFile_15 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[16]) begin
          PhysicalRegFilePlugin_logic_regFile_16 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[17]) begin
          PhysicalRegFilePlugin_logic_regFile_17 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[18]) begin
          PhysicalRegFilePlugin_logic_regFile_18 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[19]) begin
          PhysicalRegFilePlugin_logic_regFile_19 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[20]) begin
          PhysicalRegFilePlugin_logic_regFile_20 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[21]) begin
          PhysicalRegFilePlugin_logic_regFile_21 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[22]) begin
          PhysicalRegFilePlugin_logic_regFile_22 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[23]) begin
          PhysicalRegFilePlugin_logic_regFile_23 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[24]) begin
          PhysicalRegFilePlugin_logic_regFile_24 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[25]) begin
          PhysicalRegFilePlugin_logic_regFile_25 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[26]) begin
          PhysicalRegFilePlugin_logic_regFile_26 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[27]) begin
          PhysicalRegFilePlugin_logic_regFile_27 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[28]) begin
          PhysicalRegFilePlugin_logic_regFile_28 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[29]) begin
          PhysicalRegFilePlugin_logic_regFile_29 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[30]) begin
          PhysicalRegFilePlugin_logic_regFile_30 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[31]) begin
          PhysicalRegFilePlugin_logic_regFile_31 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[32]) begin
          PhysicalRegFilePlugin_logic_regFile_32 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[33]) begin
          PhysicalRegFilePlugin_logic_regFile_33 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[34]) begin
          PhysicalRegFilePlugin_logic_regFile_34 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[35]) begin
          PhysicalRegFilePlugin_logic_regFile_35 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[36]) begin
          PhysicalRegFilePlugin_logic_regFile_36 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[37]) begin
          PhysicalRegFilePlugin_logic_regFile_37 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[38]) begin
          PhysicalRegFilePlugin_logic_regFile_38 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[39]) begin
          PhysicalRegFilePlugin_logic_regFile_39 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[40]) begin
          PhysicalRegFilePlugin_logic_regFile_40 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[41]) begin
          PhysicalRegFilePlugin_logic_regFile_41 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[42]) begin
          PhysicalRegFilePlugin_logic_regFile_42 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[43]) begin
          PhysicalRegFilePlugin_logic_regFile_43 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[44]) begin
          PhysicalRegFilePlugin_logic_regFile_44 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[45]) begin
          PhysicalRegFilePlugin_logic_regFile_45 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[46]) begin
          PhysicalRegFilePlugin_logic_regFile_46 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[47]) begin
          PhysicalRegFilePlugin_logic_regFile_47 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[48]) begin
          PhysicalRegFilePlugin_logic_regFile_48 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[49]) begin
          PhysicalRegFilePlugin_logic_regFile_49 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[50]) begin
          PhysicalRegFilePlugin_logic_regFile_50 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[51]) begin
          PhysicalRegFilePlugin_logic_regFile_51 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[52]) begin
          PhysicalRegFilePlugin_logic_regFile_52 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[53]) begin
          PhysicalRegFilePlugin_logic_regFile_53 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[54]) begin
          PhysicalRegFilePlugin_logic_regFile_54 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[55]) begin
          PhysicalRegFilePlugin_logic_regFile_55 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[56]) begin
          PhysicalRegFilePlugin_logic_regFile_56 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[57]) begin
          PhysicalRegFilePlugin_logic_regFile_57 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[58]) begin
          PhysicalRegFilePlugin_logic_regFile_58 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[59]) begin
          PhysicalRegFilePlugin_logic_regFile_59 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[60]) begin
          PhysicalRegFilePlugin_logic_regFile_60 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[61]) begin
          PhysicalRegFilePlugin_logic_regFile_61 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[62]) begin
          PhysicalRegFilePlugin_logic_regFile_62 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        if(_zz_59[63]) begin
          PhysicalRegFilePlugin_logic_regFile_63 <= MulEU_MulEuPlugin_gprWritePort_data;
        end
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L134
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:134):  [normal] [PRegPlugin] Write from `MulEU.gprWritePort` to reg[%x] with data %x", MulEU_MulEuPlugin_gprWritePort_address, MulEU_MulEuPlugin_gprWritePort_data); // PhysicalRegFile.scala:L134
            end
          `endif
        `endif
      end
      if(when_PhysicalRegFile_l130_2) begin
        if(_zz_60[0]) begin
          PhysicalRegFilePlugin_logic_regFile_0 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[1]) begin
          PhysicalRegFilePlugin_logic_regFile_1 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[2]) begin
          PhysicalRegFilePlugin_logic_regFile_2 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[3]) begin
          PhysicalRegFilePlugin_logic_regFile_3 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[4]) begin
          PhysicalRegFilePlugin_logic_regFile_4 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[5]) begin
          PhysicalRegFilePlugin_logic_regFile_5 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[6]) begin
          PhysicalRegFilePlugin_logic_regFile_6 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[7]) begin
          PhysicalRegFilePlugin_logic_regFile_7 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[8]) begin
          PhysicalRegFilePlugin_logic_regFile_8 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[9]) begin
          PhysicalRegFilePlugin_logic_regFile_9 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[10]) begin
          PhysicalRegFilePlugin_logic_regFile_10 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[11]) begin
          PhysicalRegFilePlugin_logic_regFile_11 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[12]) begin
          PhysicalRegFilePlugin_logic_regFile_12 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[13]) begin
          PhysicalRegFilePlugin_logic_regFile_13 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[14]) begin
          PhysicalRegFilePlugin_logic_regFile_14 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[15]) begin
          PhysicalRegFilePlugin_logic_regFile_15 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[16]) begin
          PhysicalRegFilePlugin_logic_regFile_16 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[17]) begin
          PhysicalRegFilePlugin_logic_regFile_17 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[18]) begin
          PhysicalRegFilePlugin_logic_regFile_18 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[19]) begin
          PhysicalRegFilePlugin_logic_regFile_19 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[20]) begin
          PhysicalRegFilePlugin_logic_regFile_20 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[21]) begin
          PhysicalRegFilePlugin_logic_regFile_21 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[22]) begin
          PhysicalRegFilePlugin_logic_regFile_22 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[23]) begin
          PhysicalRegFilePlugin_logic_regFile_23 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[24]) begin
          PhysicalRegFilePlugin_logic_regFile_24 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[25]) begin
          PhysicalRegFilePlugin_logic_regFile_25 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[26]) begin
          PhysicalRegFilePlugin_logic_regFile_26 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[27]) begin
          PhysicalRegFilePlugin_logic_regFile_27 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[28]) begin
          PhysicalRegFilePlugin_logic_regFile_28 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[29]) begin
          PhysicalRegFilePlugin_logic_regFile_29 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[30]) begin
          PhysicalRegFilePlugin_logic_regFile_30 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[31]) begin
          PhysicalRegFilePlugin_logic_regFile_31 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[32]) begin
          PhysicalRegFilePlugin_logic_regFile_32 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[33]) begin
          PhysicalRegFilePlugin_logic_regFile_33 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[34]) begin
          PhysicalRegFilePlugin_logic_regFile_34 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[35]) begin
          PhysicalRegFilePlugin_logic_regFile_35 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[36]) begin
          PhysicalRegFilePlugin_logic_regFile_36 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[37]) begin
          PhysicalRegFilePlugin_logic_regFile_37 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[38]) begin
          PhysicalRegFilePlugin_logic_regFile_38 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[39]) begin
          PhysicalRegFilePlugin_logic_regFile_39 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[40]) begin
          PhysicalRegFilePlugin_logic_regFile_40 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[41]) begin
          PhysicalRegFilePlugin_logic_regFile_41 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[42]) begin
          PhysicalRegFilePlugin_logic_regFile_42 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[43]) begin
          PhysicalRegFilePlugin_logic_regFile_43 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[44]) begin
          PhysicalRegFilePlugin_logic_regFile_44 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[45]) begin
          PhysicalRegFilePlugin_logic_regFile_45 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[46]) begin
          PhysicalRegFilePlugin_logic_regFile_46 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[47]) begin
          PhysicalRegFilePlugin_logic_regFile_47 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[48]) begin
          PhysicalRegFilePlugin_logic_regFile_48 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[49]) begin
          PhysicalRegFilePlugin_logic_regFile_49 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[50]) begin
          PhysicalRegFilePlugin_logic_regFile_50 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[51]) begin
          PhysicalRegFilePlugin_logic_regFile_51 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[52]) begin
          PhysicalRegFilePlugin_logic_regFile_52 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[53]) begin
          PhysicalRegFilePlugin_logic_regFile_53 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[54]) begin
          PhysicalRegFilePlugin_logic_regFile_54 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[55]) begin
          PhysicalRegFilePlugin_logic_regFile_55 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[56]) begin
          PhysicalRegFilePlugin_logic_regFile_56 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[57]) begin
          PhysicalRegFilePlugin_logic_regFile_57 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[58]) begin
          PhysicalRegFilePlugin_logic_regFile_58 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[59]) begin
          PhysicalRegFilePlugin_logic_regFile_59 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[60]) begin
          PhysicalRegFilePlugin_logic_regFile_60 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[61]) begin
          PhysicalRegFilePlugin_logic_regFile_61 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[62]) begin
          PhysicalRegFilePlugin_logic_regFile_62 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        if(_zz_60[63]) begin
          PhysicalRegFilePlugin_logic_regFile_63 <= BranchEU_BranchEuPlugin_gprWritePort_data;
        end
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L134
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:134):  [normal] [PRegPlugin] Write from `BranchEU.gprWritePort` to reg[%x] with data %x", BranchEU_BranchEuPlugin_gprWritePort_address, BranchEU_BranchEuPlugin_gprWritePort_data); // PhysicalRegFile.scala:L134
            end
          `endif
        `endif
      end
      if(when_PhysicalRegFile_l130_3) begin
        if(_zz_61[0]) begin
          PhysicalRegFilePlugin_logic_regFile_0 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[1]) begin
          PhysicalRegFilePlugin_logic_regFile_1 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[2]) begin
          PhysicalRegFilePlugin_logic_regFile_2 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[3]) begin
          PhysicalRegFilePlugin_logic_regFile_3 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[4]) begin
          PhysicalRegFilePlugin_logic_regFile_4 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[5]) begin
          PhysicalRegFilePlugin_logic_regFile_5 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[6]) begin
          PhysicalRegFilePlugin_logic_regFile_6 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[7]) begin
          PhysicalRegFilePlugin_logic_regFile_7 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[8]) begin
          PhysicalRegFilePlugin_logic_regFile_8 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[9]) begin
          PhysicalRegFilePlugin_logic_regFile_9 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[10]) begin
          PhysicalRegFilePlugin_logic_regFile_10 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[11]) begin
          PhysicalRegFilePlugin_logic_regFile_11 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[12]) begin
          PhysicalRegFilePlugin_logic_regFile_12 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[13]) begin
          PhysicalRegFilePlugin_logic_regFile_13 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[14]) begin
          PhysicalRegFilePlugin_logic_regFile_14 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[15]) begin
          PhysicalRegFilePlugin_logic_regFile_15 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[16]) begin
          PhysicalRegFilePlugin_logic_regFile_16 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[17]) begin
          PhysicalRegFilePlugin_logic_regFile_17 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[18]) begin
          PhysicalRegFilePlugin_logic_regFile_18 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[19]) begin
          PhysicalRegFilePlugin_logic_regFile_19 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[20]) begin
          PhysicalRegFilePlugin_logic_regFile_20 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[21]) begin
          PhysicalRegFilePlugin_logic_regFile_21 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[22]) begin
          PhysicalRegFilePlugin_logic_regFile_22 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[23]) begin
          PhysicalRegFilePlugin_logic_regFile_23 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[24]) begin
          PhysicalRegFilePlugin_logic_regFile_24 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[25]) begin
          PhysicalRegFilePlugin_logic_regFile_25 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[26]) begin
          PhysicalRegFilePlugin_logic_regFile_26 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[27]) begin
          PhysicalRegFilePlugin_logic_regFile_27 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[28]) begin
          PhysicalRegFilePlugin_logic_regFile_28 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[29]) begin
          PhysicalRegFilePlugin_logic_regFile_29 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[30]) begin
          PhysicalRegFilePlugin_logic_regFile_30 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[31]) begin
          PhysicalRegFilePlugin_logic_regFile_31 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[32]) begin
          PhysicalRegFilePlugin_logic_regFile_32 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[33]) begin
          PhysicalRegFilePlugin_logic_regFile_33 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[34]) begin
          PhysicalRegFilePlugin_logic_regFile_34 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[35]) begin
          PhysicalRegFilePlugin_logic_regFile_35 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[36]) begin
          PhysicalRegFilePlugin_logic_regFile_36 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[37]) begin
          PhysicalRegFilePlugin_logic_regFile_37 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[38]) begin
          PhysicalRegFilePlugin_logic_regFile_38 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[39]) begin
          PhysicalRegFilePlugin_logic_regFile_39 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[40]) begin
          PhysicalRegFilePlugin_logic_regFile_40 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[41]) begin
          PhysicalRegFilePlugin_logic_regFile_41 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[42]) begin
          PhysicalRegFilePlugin_logic_regFile_42 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[43]) begin
          PhysicalRegFilePlugin_logic_regFile_43 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[44]) begin
          PhysicalRegFilePlugin_logic_regFile_44 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[45]) begin
          PhysicalRegFilePlugin_logic_regFile_45 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[46]) begin
          PhysicalRegFilePlugin_logic_regFile_46 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[47]) begin
          PhysicalRegFilePlugin_logic_regFile_47 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[48]) begin
          PhysicalRegFilePlugin_logic_regFile_48 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[49]) begin
          PhysicalRegFilePlugin_logic_regFile_49 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[50]) begin
          PhysicalRegFilePlugin_logic_regFile_50 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[51]) begin
          PhysicalRegFilePlugin_logic_regFile_51 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[52]) begin
          PhysicalRegFilePlugin_logic_regFile_52 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[53]) begin
          PhysicalRegFilePlugin_logic_regFile_53 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[54]) begin
          PhysicalRegFilePlugin_logic_regFile_54 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[55]) begin
          PhysicalRegFilePlugin_logic_regFile_55 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[56]) begin
          PhysicalRegFilePlugin_logic_regFile_56 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[57]) begin
          PhysicalRegFilePlugin_logic_regFile_57 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[58]) begin
          PhysicalRegFilePlugin_logic_regFile_58 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[59]) begin
          PhysicalRegFilePlugin_logic_regFile_59 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[60]) begin
          PhysicalRegFilePlugin_logic_regFile_60 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[61]) begin
          PhysicalRegFilePlugin_logic_regFile_61 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[62]) begin
          PhysicalRegFilePlugin_logic_regFile_62 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        if(_zz_61[63]) begin
          PhysicalRegFilePlugin_logic_regFile_63 <= LsuEU_LsuEuPlugin_gprWritePort_data;
        end
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L134
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:134):  [normal] [PRegPlugin] Write from `LsuEU.gprWritePort` to reg[%x] with data %x", LsuEU_LsuEuPlugin_gprWritePort_address, LsuEU_LsuEuPlugin_gprWritePort_data); // PhysicalRegFile.scala:L134
            end
          `endif
        `endif
      end
      if(when_PhysicalRegFile_l130_4) begin
        if(_zz_62[0]) begin
          PhysicalRegFilePlugin_logic_regFile_0 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[1]) begin
          PhysicalRegFilePlugin_logic_regFile_1 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[2]) begin
          PhysicalRegFilePlugin_logic_regFile_2 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[3]) begin
          PhysicalRegFilePlugin_logic_regFile_3 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[4]) begin
          PhysicalRegFilePlugin_logic_regFile_4 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[5]) begin
          PhysicalRegFilePlugin_logic_regFile_5 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[6]) begin
          PhysicalRegFilePlugin_logic_regFile_6 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[7]) begin
          PhysicalRegFilePlugin_logic_regFile_7 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[8]) begin
          PhysicalRegFilePlugin_logic_regFile_8 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[9]) begin
          PhysicalRegFilePlugin_logic_regFile_9 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[10]) begin
          PhysicalRegFilePlugin_logic_regFile_10 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[11]) begin
          PhysicalRegFilePlugin_logic_regFile_11 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[12]) begin
          PhysicalRegFilePlugin_logic_regFile_12 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[13]) begin
          PhysicalRegFilePlugin_logic_regFile_13 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[14]) begin
          PhysicalRegFilePlugin_logic_regFile_14 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[15]) begin
          PhysicalRegFilePlugin_logic_regFile_15 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[16]) begin
          PhysicalRegFilePlugin_logic_regFile_16 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[17]) begin
          PhysicalRegFilePlugin_logic_regFile_17 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[18]) begin
          PhysicalRegFilePlugin_logic_regFile_18 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[19]) begin
          PhysicalRegFilePlugin_logic_regFile_19 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[20]) begin
          PhysicalRegFilePlugin_logic_regFile_20 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[21]) begin
          PhysicalRegFilePlugin_logic_regFile_21 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[22]) begin
          PhysicalRegFilePlugin_logic_regFile_22 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[23]) begin
          PhysicalRegFilePlugin_logic_regFile_23 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[24]) begin
          PhysicalRegFilePlugin_logic_regFile_24 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[25]) begin
          PhysicalRegFilePlugin_logic_regFile_25 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[26]) begin
          PhysicalRegFilePlugin_logic_regFile_26 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[27]) begin
          PhysicalRegFilePlugin_logic_regFile_27 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[28]) begin
          PhysicalRegFilePlugin_logic_regFile_28 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[29]) begin
          PhysicalRegFilePlugin_logic_regFile_29 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[30]) begin
          PhysicalRegFilePlugin_logic_regFile_30 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[31]) begin
          PhysicalRegFilePlugin_logic_regFile_31 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[32]) begin
          PhysicalRegFilePlugin_logic_regFile_32 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[33]) begin
          PhysicalRegFilePlugin_logic_regFile_33 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[34]) begin
          PhysicalRegFilePlugin_logic_regFile_34 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[35]) begin
          PhysicalRegFilePlugin_logic_regFile_35 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[36]) begin
          PhysicalRegFilePlugin_logic_regFile_36 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[37]) begin
          PhysicalRegFilePlugin_logic_regFile_37 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[38]) begin
          PhysicalRegFilePlugin_logic_regFile_38 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[39]) begin
          PhysicalRegFilePlugin_logic_regFile_39 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[40]) begin
          PhysicalRegFilePlugin_logic_regFile_40 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[41]) begin
          PhysicalRegFilePlugin_logic_regFile_41 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[42]) begin
          PhysicalRegFilePlugin_logic_regFile_42 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[43]) begin
          PhysicalRegFilePlugin_logic_regFile_43 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[44]) begin
          PhysicalRegFilePlugin_logic_regFile_44 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[45]) begin
          PhysicalRegFilePlugin_logic_regFile_45 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[46]) begin
          PhysicalRegFilePlugin_logic_regFile_46 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[47]) begin
          PhysicalRegFilePlugin_logic_regFile_47 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[48]) begin
          PhysicalRegFilePlugin_logic_regFile_48 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[49]) begin
          PhysicalRegFilePlugin_logic_regFile_49 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[50]) begin
          PhysicalRegFilePlugin_logic_regFile_50 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[51]) begin
          PhysicalRegFilePlugin_logic_regFile_51 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[52]) begin
          PhysicalRegFilePlugin_logic_regFile_52 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[53]) begin
          PhysicalRegFilePlugin_logic_regFile_53 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[54]) begin
          PhysicalRegFilePlugin_logic_regFile_54 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[55]) begin
          PhysicalRegFilePlugin_logic_regFile_55 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[56]) begin
          PhysicalRegFilePlugin_logic_regFile_56 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[57]) begin
          PhysicalRegFilePlugin_logic_regFile_57 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[58]) begin
          PhysicalRegFilePlugin_logic_regFile_58 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[59]) begin
          PhysicalRegFilePlugin_logic_regFile_59 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[60]) begin
          PhysicalRegFilePlugin_logic_regFile_60 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[61]) begin
          PhysicalRegFilePlugin_logic_regFile_61 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[62]) begin
          PhysicalRegFilePlugin_logic_regFile_62 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        if(_zz_62[63]) begin
          PhysicalRegFilePlugin_logic_regFile_63 <= LoadQueuePlugin_hw_prfWritePort_data;
        end
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // PhysicalRegFile.scala:L134
          `else
            if(!1'b0) begin
              $display("NOTE(PhysicalRegFile.scala:134):  [normal] [PRegPlugin] Write from `LQ.gprWritePort` to reg[%x] with data %x", LoadQueuePlugin_hw_prfWritePort_address, LoadQueuePlugin_hw_prfWritePort_data); // PhysicalRegFile.scala:L134
            end
          `endif
        `endif
      end
      StoreBufferPlugin_logic_registeredFlush_valid <= StoreBufferPlugin_logic_flushInProgress;
      StoreBufferPlugin_logic_registeredFlush_targetRobPtr <= ROBPlugin_aggregatedFlushSignal_payload_targetRobPtr;
      if(when_StoreBufferPlugin_l316) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L317
          `else
            if(!1'b0) begin
              $display("FAILURE Got isIO but no MMIO service."); // StoreBufferPlugin.scala:L317
              $finish;
            end
          `endif
        `endif
      end
      if(StoreBufferPlugin_logic_mmioCmdFired) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L408
          `else
            if(!1'b0) begin
              $display("NOTE(StoreBufferPlugin.scala:408):  [SQ] CMD_FIRED_MMIO: robPtr=%x (slotIdx=0), addr=%x", StoreBufferPlugin_logic_slots_0_robPtr, StoreBufferPlugin_logic_slots_0_addr); // StoreBufferPlugin.scala:L408
            end
          `endif
        `endif
      end
      if(StoreBufferPlugin_logic_mmioResponseForHead) begin
        if(CoreMemSysPlugin_logic_writeBridges_0_io_gmbIn_write_rsp_payload_error) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // StoreBufferPlugin.scala:L440
            `else
              if(!1'b0) begin
                $display("NOTE(StoreBufferPlugin.scala:440):  [SQ-MMIO] MMIO RSP_ERROR received for robPtr=%x.", StoreBufferPlugin_logic_slots_0_robPtr); // StoreBufferPlugin.scala:L440
              end
            `endif
          `endif
        end else begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // StoreBufferPlugin.scala:L445
            `else
              if(!1'b0) begin
                $display("NOTE(StoreBufferPlugin.scala:445):  [SQ-MMIO] MMIO RSP_SUCCESS received for robPtr=%x.", StoreBufferPlugin_logic_slots_0_robPtr); // StoreBufferPlugin.scala:L445
              end
            `endif
          `endif
        end
      end
      if(oneShot_25_io_pulseOut) begin
        if(when_Debug_l71_11) begin
          _zz_when_Debug_l71 <= {2'd0, _zz_when_Debug_l71_12};
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // Debug.scala:L73
            `else
              if(!1'b0) begin
                $display("NOTE(Debug.scala:73):  [DbgSvc] Set (expect incremental) value to 0x%x", _zz_when_Debug_l71_12); // Debug.scala:L73
              end
            `endif
          `endif
        end
      end
      if(when_StoreBufferPlugin_l498) begin
        if(when_StoreBufferPlugin_l504) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // StoreBufferPlugin.scala:L507
            `else
              if(!1'b0) begin
                $display("NOTE(StoreBufferPlugin.scala:507):  [SQ] COMMIT_DETECT: robPtr=%x (slotIdx=0) will be marked as committed next cycle.", StoreBufferPlugin_logic_slots_0_robPtr); // StoreBufferPlugin.scala:L507
              end
            `endif
          `endif
        end
      end
      if(when_StoreBufferPlugin_l498_1) begin
        if(when_StoreBufferPlugin_l504_1) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // StoreBufferPlugin.scala:L507
            `else
              if(!1'b0) begin
                $display("NOTE(StoreBufferPlugin.scala:507):  [SQ] COMMIT_DETECT: robPtr=%x (slotIdx=1) will be marked as committed next cycle.", StoreBufferPlugin_logic_slots_1_robPtr); // StoreBufferPlugin.scala:L507
              end
            `endif
          `endif
        end
      end
      if(when_StoreBufferPlugin_l498_2) begin
        if(when_StoreBufferPlugin_l504_2) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // StoreBufferPlugin.scala:L507
            `else
              if(!1'b0) begin
                $display("NOTE(StoreBufferPlugin.scala:507):  [SQ] COMMIT_DETECT: robPtr=%x (slotIdx=2) will be marked as committed next cycle.", StoreBufferPlugin_logic_slots_2_robPtr); // StoreBufferPlugin.scala:L507
              end
            `endif
          `endif
        end
      end
      if(when_StoreBufferPlugin_l498_3) begin
        if(when_StoreBufferPlugin_l504_3) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // StoreBufferPlugin.scala:L507
            `else
              if(!1'b0) begin
                $display("NOTE(StoreBufferPlugin.scala:507):  [SQ] COMMIT_DETECT: robPtr=%x (slotIdx=3) will be marked as committed next cycle.", StoreBufferPlugin_logic_slots_3_robPtr); // StoreBufferPlugin.scala:L507
              end
            `endif
          `endif
        end
      end
      StoreBufferPlugin_logic_registeredCommitUpdate_validMask <= StoreBufferPlugin_logic_commitUpdateInfo_validMask;
      if(when_StoreBufferPlugin_l525) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L528
          `else
            if(!1'b0) begin
              $display("NOTE(StoreBufferPlugin.scala:528):  [SQ] FLUSH (Exec): Invalidating slotIdx=0 (robPtr=%x) by ROB flush.", StoreBufferPlugin_logic_slots_0_robPtr); // StoreBufferPlugin.scala:L528
            end
          `endif
        `endif
      end
      if(when_StoreBufferPlugin_l525_1) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L528
          `else
            if(!1'b0) begin
              $display("NOTE(StoreBufferPlugin.scala:528):  [SQ] FLUSH (Exec): Invalidating slotIdx=1 (robPtr=%x) by ROB flush.", StoreBufferPlugin_logic_slots_1_robPtr); // StoreBufferPlugin.scala:L528
            end
          `endif
        `endif
      end
      if(when_StoreBufferPlugin_l525_2) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L528
          `else
            if(!1'b0) begin
              $display("NOTE(StoreBufferPlugin.scala:528):  [SQ] FLUSH (Exec): Invalidating slotIdx=2 (robPtr=%x) by ROB flush.", StoreBufferPlugin_logic_slots_2_robPtr); // StoreBufferPlugin.scala:L528
            end
          `endif
        `endif
      end
      if(when_StoreBufferPlugin_l525_3) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L528
          `else
            if(!1'b0) begin
              $display("NOTE(StoreBufferPlugin.scala:528):  [SQ] FLUSH (Exec): Invalidating slotIdx=3 (robPtr=%x) by ROB flush.", StoreBufferPlugin_logic_slots_3_robPtr); // StoreBufferPlugin.scala:L528
            end
          `endif
        `endif
      end
      if(when_StoreBufferPlugin_l555) begin
        if(StoreBufferPlugin_logic_slotsAfterUpdates_0_isFlush) begin
          if(StoreBufferPlugin_logic_operationDone) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // StoreBufferPlugin.scala:L560
              `else
                if(!1'b0) begin
                  $display("NOTE(StoreBufferPlugin.scala:560):  [SQ] POP_FLUSH: robPtr=%x", StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr); // StoreBufferPlugin.scala:L560
                end
              `endif
            `endif
          end
        end else begin
          if(StoreBufferPlugin_logic_slotsAfterUpdates_0_hasEarlyException) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // StoreBufferPlugin.scala:L567
              `else
                if(!1'b0) begin
                  $display("NOTE(StoreBufferPlugin.scala:567):  [SQ] POP_EARLY_EXCEPTION: robPtr=%x", StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr); // StoreBufferPlugin.scala:L567
                end
              `endif
            `endif
          end else begin
            if(StoreBufferPlugin_logic_operationDone) begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // StoreBufferPlugin.scala:L572
                `else
                  if(!1'b0) begin
                    $display("NOTE(StoreBufferPlugin.scala:572):  [SQ] POP_NORMAL_STORE/MMIO: robPtr=%x, isIO=%x", StoreBufferPlugin_logic_slotsAfterUpdates_0_robPtr, StoreBufferPlugin_logic_slotsAfterUpdates_0_isIO); // StoreBufferPlugin.scala:L572
                  end
                `endif
              `endif
            end
          end
        end
      end
      if(StoreBufferPlugin_hw_sqQueryPort_cmd_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L613
          `else
            if(!1'b0) begin
              $display("NOTE(StoreBufferPlugin.scala:613):  [SQ-Fwd] Query: valid=%x robPtr=%x addr=%x size=%s", StoreBufferPlugin_hw_sqQueryPort_cmd_valid, StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr, StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address, StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size_string); // StoreBufferPlugin.scala:L613
            end
          `endif
        `endif
      end
      if(when_StoreBufferPlugin_l672) begin
        if(when_StoreBufferPlugin_l678) begin
          if(when_StoreBufferPlugin_l681) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // StoreBufferPlugin.scala:L682
              `else
                if(!1'b0) begin
                  $display("NOTE(StoreBufferPlugin.scala:682):  [SQ-Fwd] STALL_DATA_NOT_READY (Slot Status): slot=%x (LoadAddr=%x, StoreAddr=%x)reason: waitRsp=%x, isWaitingForRefill=%x, isWaitingForWb=%x", StoreBufferPlugin_logic_slots_0_robPtr, _zz_when_StoreBufferPlugin_l678_4, _zz_when_StoreBufferPlugin_l678_5, StoreBufferPlugin_logic_slots_0_waitRsp, StoreBufferPlugin_logic_slots_0_isWaitingForRefill, StoreBufferPlugin_logic_slots_0_isWaitingForWb); // StoreBufferPlugin.scala:L682
                end
              `endif
            `endif
          end
        end
      end
      if(when_StoreBufferPlugin_l672_1) begin
        if(when_StoreBufferPlugin_l678_1) begin
          if(when_StoreBufferPlugin_l681_1) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // StoreBufferPlugin.scala:L682
              `else
                if(!1'b0) begin
                  $display("NOTE(StoreBufferPlugin.scala:682):  [SQ-Fwd] STALL_DATA_NOT_READY (Slot Status): slot=%x (LoadAddr=%x, StoreAddr=%x)reason: waitRsp=%x, isWaitingForRefill=%x, isWaitingForWb=%x", StoreBufferPlugin_logic_slots_1_robPtr, _zz_when_StoreBufferPlugin_l678_10, _zz_when_StoreBufferPlugin_l678_11, StoreBufferPlugin_logic_slots_1_waitRsp, StoreBufferPlugin_logic_slots_1_isWaitingForRefill, StoreBufferPlugin_logic_slots_1_isWaitingForWb); // StoreBufferPlugin.scala:L682
                end
              `endif
            `endif
          end
        end
      end
      if(when_StoreBufferPlugin_l672_2) begin
        if(when_StoreBufferPlugin_l678_2) begin
          if(when_StoreBufferPlugin_l681_2) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // StoreBufferPlugin.scala:L682
              `else
                if(!1'b0) begin
                  $display("NOTE(StoreBufferPlugin.scala:682):  [SQ-Fwd] STALL_DATA_NOT_READY (Slot Status): slot=%x (LoadAddr=%x, StoreAddr=%x)reason: waitRsp=%x, isWaitingForRefill=%x, isWaitingForWb=%x", StoreBufferPlugin_logic_slots_2_robPtr, _zz_when_StoreBufferPlugin_l678_16, _zz_when_StoreBufferPlugin_l678_17, StoreBufferPlugin_logic_slots_2_waitRsp, StoreBufferPlugin_logic_slots_2_isWaitingForRefill, StoreBufferPlugin_logic_slots_2_isWaitingForWb); // StoreBufferPlugin.scala:L682
                end
              `endif
            `endif
          end
        end
      end
      if(when_StoreBufferPlugin_l672_3) begin
        if(when_StoreBufferPlugin_l678_3) begin
          if(when_StoreBufferPlugin_l681_3) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // StoreBufferPlugin.scala:L682
              `else
                if(!1'b0) begin
                  $display("NOTE(StoreBufferPlugin.scala:682):  [SQ-Fwd] STALL_DATA_NOT_READY (Slot Status): slot=%x (LoadAddr=%x, StoreAddr=%x)reason: waitRsp=%x, isWaitingForRefill=%x, isWaitingForWb=%x", StoreBufferPlugin_logic_slots_3_robPtr, _zz_when_StoreBufferPlugin_l678_22, _zz_when_StoreBufferPlugin_l678_23, StoreBufferPlugin_logic_slots_3_waitRsp, StoreBufferPlugin_logic_slots_3_isWaitingForRefill, StoreBufferPlugin_logic_slots_3_isWaitingForWb); // StoreBufferPlugin.scala:L682
                end
              `endif
            `endif
          end
        end
      end
      if(StoreBufferPlugin_hw_sqQueryPort_cmd_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L711
          `else
            if(!1'b0) begin
              $display("NOTE(StoreBufferPlugin.scala:711):  [SQ-Fwd] Query: SqQuery(robPtr=%x,address=%x,size=%s)", StoreBufferPlugin_hw_sqQueryPort_cmd_payload_robPtr, StoreBufferPlugin_hw_sqQueryPort_cmd_payload_address, StoreBufferPlugin_hw_sqQueryPort_cmd_payload_size_string); // StoreBufferPlugin.scala:L711
            end
          `endif
        `endif
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // StoreBufferPlugin.scala:L712
          `else
            if(!1'b0) begin
              $display("NOTE(StoreBufferPlugin.scala:712):  [SQ-Fwd] Rsp: SqQueryRsp(hit=%x,data=%x,olderStoreHasUnknownAddress=%x,olderStoreDataNotReady=%x)", StoreBufferPlugin_hw_sqQueryPort_rsp_hit, StoreBufferPlugin_hw_sqQueryPort_rsp_data, StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreHasUnknownAddress, StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreDataNotReady); // StoreBufferPlugin.scala:L712
            end
          `endif
        `endif
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // StoreBufferPlugin.scala:L714
        `else
          if(!1'b0) begin
            $display("NOTE(StoreBufferPlugin.scala:714):  [SQ-Fwd] Result: hitMask=%x (loadMask=%x), allHit=%x, finalRsp.hit=%x", StoreBufferPlugin_logic_forwardingLogic_forwardingResult_hitMask, StoreBufferPlugin_logic_forwardingLogic_loadMask, StoreBufferPlugin_logic_forwardingLogic_allRequiredBytesHit, StoreBufferPlugin_hw_sqQueryPort_rsp_hit); // StoreBufferPlugin.scala:L714
          end
        `endif
      `endif
      StoreBufferPlugin_logic_slots_0_isFlush <= StoreBufferPlugin_logic_slotsNext_0_isFlush;
      StoreBufferPlugin_logic_slots_0_addr <= StoreBufferPlugin_logic_slotsNext_0_addr;
      StoreBufferPlugin_logic_slots_0_data <= StoreBufferPlugin_logic_slotsNext_0_data;
      StoreBufferPlugin_logic_slots_0_be <= StoreBufferPlugin_logic_slotsNext_0_be;
      StoreBufferPlugin_logic_slots_0_robPtr <= StoreBufferPlugin_logic_slotsNext_0_robPtr;
      StoreBufferPlugin_logic_slots_0_accessSize <= StoreBufferPlugin_logic_slotsNext_0_accessSize;
      StoreBufferPlugin_logic_slots_0_isIO <= StoreBufferPlugin_logic_slotsNext_0_isIO;
      StoreBufferPlugin_logic_slots_0_valid <= StoreBufferPlugin_logic_slotsNext_0_valid;
      StoreBufferPlugin_logic_slots_0_hasEarlyException <= StoreBufferPlugin_logic_slotsNext_0_hasEarlyException;
      StoreBufferPlugin_logic_slots_0_earlyExceptionCode <= StoreBufferPlugin_logic_slotsNext_0_earlyExceptionCode;
      StoreBufferPlugin_logic_slots_0_isCommitted <= StoreBufferPlugin_logic_slotsNext_0_isCommitted;
      StoreBufferPlugin_logic_slots_0_sentCmd <= StoreBufferPlugin_logic_slotsNext_0_sentCmd;
      StoreBufferPlugin_logic_slots_0_waitRsp <= StoreBufferPlugin_logic_slotsNext_0_waitRsp;
      StoreBufferPlugin_logic_slots_0_isWaitingForRefill <= StoreBufferPlugin_logic_slotsNext_0_isWaitingForRefill;
      StoreBufferPlugin_logic_slots_0_isWaitingForWb <= StoreBufferPlugin_logic_slotsNext_0_isWaitingForWb;
      StoreBufferPlugin_logic_slots_0_refillSlotToWatch <= StoreBufferPlugin_logic_slotsNext_0_refillSlotToWatch;
      StoreBufferPlugin_logic_slots_1_isFlush <= StoreBufferPlugin_logic_slotsNext_1_isFlush;
      StoreBufferPlugin_logic_slots_1_addr <= StoreBufferPlugin_logic_slotsNext_1_addr;
      StoreBufferPlugin_logic_slots_1_data <= StoreBufferPlugin_logic_slotsNext_1_data;
      StoreBufferPlugin_logic_slots_1_be <= StoreBufferPlugin_logic_slotsNext_1_be;
      StoreBufferPlugin_logic_slots_1_robPtr <= StoreBufferPlugin_logic_slotsNext_1_robPtr;
      StoreBufferPlugin_logic_slots_1_accessSize <= StoreBufferPlugin_logic_slotsNext_1_accessSize;
      StoreBufferPlugin_logic_slots_1_isIO <= StoreBufferPlugin_logic_slotsNext_1_isIO;
      StoreBufferPlugin_logic_slots_1_valid <= StoreBufferPlugin_logic_slotsNext_1_valid;
      StoreBufferPlugin_logic_slots_1_hasEarlyException <= StoreBufferPlugin_logic_slotsNext_1_hasEarlyException;
      StoreBufferPlugin_logic_slots_1_earlyExceptionCode <= StoreBufferPlugin_logic_slotsNext_1_earlyExceptionCode;
      StoreBufferPlugin_logic_slots_1_isCommitted <= StoreBufferPlugin_logic_slotsNext_1_isCommitted;
      StoreBufferPlugin_logic_slots_1_sentCmd <= StoreBufferPlugin_logic_slotsNext_1_sentCmd;
      StoreBufferPlugin_logic_slots_1_waitRsp <= StoreBufferPlugin_logic_slotsNext_1_waitRsp;
      StoreBufferPlugin_logic_slots_1_isWaitingForRefill <= StoreBufferPlugin_logic_slotsNext_1_isWaitingForRefill;
      StoreBufferPlugin_logic_slots_1_isWaitingForWb <= StoreBufferPlugin_logic_slotsNext_1_isWaitingForWb;
      StoreBufferPlugin_logic_slots_1_refillSlotToWatch <= StoreBufferPlugin_logic_slotsNext_1_refillSlotToWatch;
      StoreBufferPlugin_logic_slots_2_isFlush <= StoreBufferPlugin_logic_slotsNext_2_isFlush;
      StoreBufferPlugin_logic_slots_2_addr <= StoreBufferPlugin_logic_slotsNext_2_addr;
      StoreBufferPlugin_logic_slots_2_data <= StoreBufferPlugin_logic_slotsNext_2_data;
      StoreBufferPlugin_logic_slots_2_be <= StoreBufferPlugin_logic_slotsNext_2_be;
      StoreBufferPlugin_logic_slots_2_robPtr <= StoreBufferPlugin_logic_slotsNext_2_robPtr;
      StoreBufferPlugin_logic_slots_2_accessSize <= StoreBufferPlugin_logic_slotsNext_2_accessSize;
      StoreBufferPlugin_logic_slots_2_isIO <= StoreBufferPlugin_logic_slotsNext_2_isIO;
      StoreBufferPlugin_logic_slots_2_valid <= StoreBufferPlugin_logic_slotsNext_2_valid;
      StoreBufferPlugin_logic_slots_2_hasEarlyException <= StoreBufferPlugin_logic_slotsNext_2_hasEarlyException;
      StoreBufferPlugin_logic_slots_2_earlyExceptionCode <= StoreBufferPlugin_logic_slotsNext_2_earlyExceptionCode;
      StoreBufferPlugin_logic_slots_2_isCommitted <= StoreBufferPlugin_logic_slotsNext_2_isCommitted;
      StoreBufferPlugin_logic_slots_2_sentCmd <= StoreBufferPlugin_logic_slotsNext_2_sentCmd;
      StoreBufferPlugin_logic_slots_2_waitRsp <= StoreBufferPlugin_logic_slotsNext_2_waitRsp;
      StoreBufferPlugin_logic_slots_2_isWaitingForRefill <= StoreBufferPlugin_logic_slotsNext_2_isWaitingForRefill;
      StoreBufferPlugin_logic_slots_2_isWaitingForWb <= StoreBufferPlugin_logic_slotsNext_2_isWaitingForWb;
      StoreBufferPlugin_logic_slots_2_refillSlotToWatch <= StoreBufferPlugin_logic_slotsNext_2_refillSlotToWatch;
      StoreBufferPlugin_logic_slots_3_isFlush <= StoreBufferPlugin_logic_slotsNext_3_isFlush;
      StoreBufferPlugin_logic_slots_3_addr <= StoreBufferPlugin_logic_slotsNext_3_addr;
      StoreBufferPlugin_logic_slots_3_data <= StoreBufferPlugin_logic_slotsNext_3_data;
      StoreBufferPlugin_logic_slots_3_be <= StoreBufferPlugin_logic_slotsNext_3_be;
      StoreBufferPlugin_logic_slots_3_robPtr <= StoreBufferPlugin_logic_slotsNext_3_robPtr;
      StoreBufferPlugin_logic_slots_3_accessSize <= StoreBufferPlugin_logic_slotsNext_3_accessSize;
      StoreBufferPlugin_logic_slots_3_isIO <= StoreBufferPlugin_logic_slotsNext_3_isIO;
      StoreBufferPlugin_logic_slots_3_valid <= StoreBufferPlugin_logic_slotsNext_3_valid;
      StoreBufferPlugin_logic_slots_3_hasEarlyException <= StoreBufferPlugin_logic_slotsNext_3_hasEarlyException;
      StoreBufferPlugin_logic_slots_3_earlyExceptionCode <= StoreBufferPlugin_logic_slotsNext_3_earlyExceptionCode;
      StoreBufferPlugin_logic_slots_3_isCommitted <= StoreBufferPlugin_logic_slotsNext_3_isCommitted;
      StoreBufferPlugin_logic_slots_3_sentCmd <= StoreBufferPlugin_logic_slotsNext_3_sentCmd;
      StoreBufferPlugin_logic_slots_3_waitRsp <= StoreBufferPlugin_logic_slotsNext_3_waitRsp;
      StoreBufferPlugin_logic_slots_3_isWaitingForRefill <= StoreBufferPlugin_logic_slotsNext_3_isWaitingForRefill;
      StoreBufferPlugin_logic_slots_3_isWaitingForWb <= StoreBufferPlugin_logic_slotsNext_3_isWaitingForWb;
      StoreBufferPlugin_logic_slots_3_refillSlotToWatch <= StoreBufferPlugin_logic_slotsNext_3_refillSlotToWatch;
      if(LinkerPlugin_logic_allWakeupFlows_0_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // WakeupPlugin.scala:L75
          `else
            if(!1'b0) begin
              $display("NOTE(WakeupPlugin.scala:75):  [normal] WakeupPlugin: Broadcasting from source[0] for physReg=%x", LinkerPlugin_logic_allWakeupFlows_0_payload_physRegIdx); // WakeupPlugin.scala:L75
            end
          `endif
        `endif
      end
      if(LinkerPlugin_logic_allWakeupFlows_1_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // WakeupPlugin.scala:L75
          `else
            if(!1'b0) begin
              $display("NOTE(WakeupPlugin.scala:75):  [normal] WakeupPlugin: Broadcasting from source[1] for physReg=%x", LinkerPlugin_logic_allWakeupFlows_1_payload_physRegIdx); // WakeupPlugin.scala:L75
            end
          `endif
        `endif
      end
      if(LinkerPlugin_logic_allWakeupFlows_2_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // WakeupPlugin.scala:L75
          `else
            if(!1'b0) begin
              $display("NOTE(WakeupPlugin.scala:75):  [normal] WakeupPlugin: Broadcasting from source[2] for physReg=%x", LinkerPlugin_logic_allWakeupFlows_2_payload_physRegIdx); // WakeupPlugin.scala:L75
            end
          `endif
        `endif
      end
      if(LinkerPlugin_logic_allWakeupFlows_3_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // WakeupPlugin.scala:L75
          `else
            if(!1'b0) begin
              $display("NOTE(WakeupPlugin.scala:75):  [normal] WakeupPlugin: Broadcasting from source[3] for physReg=%x", LinkerPlugin_logic_allWakeupFlows_3_payload_physRegIdx); // WakeupPlugin.scala:L75
            end
          `endif
        `endif
      end
      if(LinkerPlugin_logic_allWakeupFlows_4_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // WakeupPlugin.scala:L75
          `else
            if(!1'b0) begin
              $display("NOTE(WakeupPlugin.scala:75):  [normal] WakeupPlugin: Broadcasting from source[4] for physReg=%x", LinkerPlugin_logic_allWakeupFlows_4_payload_physRegIdx); // WakeupPlugin.scala:L75
            end
          `endif
        `endif
      end
      if(CheckpointManagerPlugin_setup_btRestorePort_valid) begin
        BusyTablePlugin_early_setup_busyTableReg <= CheckpointManagerPlugin_setup_btRestorePort_payload_busyBits;
      end else begin
        BusyTablePlugin_early_setup_busyTableReg <= BusyTablePlugin_logic_busyTableNext;
      end
      FetchPipelinePlugin_logic_retryIdCounter_value <= FetchPipelinePlugin_logic_retryIdCounter_valueNext;
      if(FetchPipelinePlugin_logic_dispatcher_io_softRedirect_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L244
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:244):  [notice] [33m[%x] !!!!GOT A SOFT REDIRECT to 0x%x!!!![0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_dispatcher_io_softRedirect_payload); // FetchPipelinePlugin2.scala:L244
            end
          `endif
        `endif
      end
      if(FetchPipelinePlugin_logic_hardRedirect_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L264
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:264):  [notice] [33m[%x] !!!!GOT A HARD FLUSH to %x[0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_hardRedirect_payload); // FetchPipelinePlugin2.scala:L264
            end
          `endif
        `endif
      end
      if(FetchPipelinePlugin_logic_dispatcher_io_softRedirect_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L267
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:267):  [notice] [33m[%x] !!!!GOT A SOFT FLUSH to %x[0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_dispatcher_io_softRedirect_payload); // FetchPipelinePlugin2.scala:L267
            end
          `endif
        `endif
      end
      if(io_pop_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L273
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:273):  [notice] [33m[%x] output a instr to decoder: PC=0x%x, instr=0x%x[0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_pc, FetchPipelinePlugin_setup_fetchOutput_io_pop_payload_instruction); // FetchPipelinePlugin2.scala:L273
            end
          `endif
        `endif
      end
      FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value <= FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_valueNext;
      if(FetchPipelinePlugin_logic_doAnyFlush) begin
        FetchPipelinePlugin_logic_isDrainingCacheRspReg <= 1'b1;
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L286
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:286):  [notice] [33m[%x] Draining the pipeline due to a flush. iCacheInFlightToDrainCounter.value=%x[0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value); // FetchPipelinePlugin2.scala:L286
            end
          `endif
        `endif
      end
      if(FetchPipelinePlugin_logic_isDrainingCacheRspReg) begin
        if(when_FetchPipelinePlugin2_l289) begin
          FetchPipelinePlugin_logic_isDrainingCacheRspReg <= 1'b0;
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // FetchPipelinePlugin2.scala:L291
            `else
              if(!1'b0) begin
                $display("NOTE(FetchPipelinePlugin2.scala:291):  [success] [32m[%x] Pipeline still has %x cycles to drain[0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value); // FetchPipelinePlugin2.scala:L291
              end
            `endif
          `endif
        end else begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // FetchPipelinePlugin2.scala:L294
            `else
              if(!1'b0) begin
                $display("NOTE(FetchPipelinePlugin2.scala:294):  [notice] [33m[%x] Pipeline still has %x cycles to drain[0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value); // FetchPipelinePlugin2.scala:L294
              end
            `endif
          `endif
        end
      end
      if(FetchPipelinePlugin_logic_hardRedirect_valid) begin
        FetchPipelinePlugin_logic_s1_logic_fetchPcReg <= FetchPipelinePlugin_logic_hardRedirect_payload;
        FetchPipelinePlugin_logic_retryCmd_lock <= 1'b0;
        FetchPipelinePlugin_logic_s1_logic_lastRetryIdReg <= 2'b00;
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L346
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:346):  [normal] [%x] FETCH-S1: fetchPcReg reset to %x due to hard flush, retry cancelled.", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_hardRedirect_payload); // FetchPipelinePlugin2.scala:L346
            end
          `endif
        `endif
      end else begin
        if(FetchPipelinePlugin_logic_dispatcher_io_softRedirect_valid) begin
          FetchPipelinePlugin_logic_s1_logic_fetchPcReg <= FetchPipelinePlugin_logic_dispatcher_io_softRedirect_payload;
          FetchPipelinePlugin_logic_retryCmd_lock <= 1'b0;
          FetchPipelinePlugin_logic_s1_logic_lastRetryIdReg <= 2'b00;
        end else begin
          if(FetchPipelinePlugin_logic_s1_logic_needRedo) begin
            FetchPipelinePlugin_logic_s1_logic_fetchPcReg <= _zz_FetchPipelinePlugin_logic_s1_logic_fetchPcReg;
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // FetchPipelinePlugin2.scala:L359
              `else
                if(!1'b0) begin
                  $display("NOTE(FetchPipelinePlugin2.scala:359):  [normal] [%x] FETCH-S1: Correcting fetchPcReg for next cycle to 0x%x", FetchPipelinePlugin_dbg_cycles, _zz_FetchPipelinePlugin_logic_s1_logic_fetchPcReg); // FetchPipelinePlugin2.scala:L359
                end
              `endif
            `endif
          end else begin
            if(when_FetchPipelinePlugin2_l361) begin
              FetchPipelinePlugin_logic_s1_logic_fetchPcReg <= FetchPipelinePlugin_logic_s1_logic_nextLinePc;
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // FetchPipelinePlugin2.scala:L363
                `else
                  if(!1'b0) begin
                    $display("NOTE(FetchPipelinePlugin2.scala:363):  [normal] [%x] FETCH-S1: fetchPcReg updated to %x (from raw PC=0x%x)", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_s1_logic_nextLinePc, s1_PC_Gen_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC); // FetchPipelinePlugin2.scala:L363
                  end
                `endif
              `endif
            end
          end
        end
      end
      if(when_FetchPipelinePlugin2_l367) begin
        FetchPipelinePlugin_logic_s1_logic_lastRetryIdReg <= FetchPipelinePlugin_logic_retryCmd_id;
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L369
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:369):  [notice] [33m[%x] FETCH-S1: Acting on retry for ID %x, PC=0x%x. Locking this ID in s1.[0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_retryCmd_id, FetchPipelinePlugin_logic_retryCmd_pc); // FetchPipelinePlugin2.scala:L369
            end
          `endif
        `endif
      end
      if(when_FetchPipelinePlugin2_l380) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L382
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:382):  [normal] [%x] FETCH-S1: Halting due to isDrainingCacheRspReg=%x, fetchDisabled=%x, iCacheInFlightToDrainCounter.value=%xretryCmd.lock=%x retryCmd.id=%x === lastRetryIdReg=%x", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_isDrainingCacheRspReg, FetchPipelinePlugin_logic_s1_logic_fetchDisabled, FetchPipelinePlugin_logic_iCacheInFlightToDrainCounter_value, FetchPipelinePlugin_logic_retryCmd_lock, FetchPipelinePlugin_logic_retryCmd_id, FetchPipelinePlugin_logic_s1_logic_lastRetryIdReg); // FetchPipelinePlugin2.scala:L382
            end
          `endif
        `endif
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // FetchPipelinePlugin2.scala:L434
        `else
          if(!1'b0) begin
            $display("NOTE(FetchPipelinePlugin2.scala:434):  [normal] [%x] FETCH-S4: Handling Rsp for PC=0x%x? %x because isFiring=%x, iCacheRsp.valid=%x, isDrainingCacheRspReg=%x", FetchPipelinePlugin_dbg_cycles, s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC, FetchPipelinePlugin_logic_s4_logic_handleRsp, s4_Predecode_isFiring, ICachePlugin_port_rsp_valid, FetchPipelinePlugin_logic_isDrainingCacheRspReg); // FetchPipelinePlugin2.scala:L434
          end
        `endif
      `endif
      if(FetchPipelinePlugin_logic_s4_logic_backpressureRedo) begin
        if(when_FetchPipelinePlugin2_l442) begin
          FetchPipelinePlugin_logic_retryCmd_lock <= 1'b1;
          FetchPipelinePlugin_logic_retryCmd_pc <= s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC;
          FetchPipelinePlugin_logic_retryCmd_id <= FetchPipelinePlugin_logic_retryIdCounter_value;
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // FetchPipelinePlugin2.scala:L448
            `else
              if(!1'b0) begin
                $display("NOTE(FetchPipelinePlugin2.scala:448):  [notice] [33m[FETCH-S4] BACKPRESSURE REDO requested for raw PC=0x%x, ID=%x because downstream FIFO is full, retryCmd.id=%x.[0m", s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC, ICachePlugin_port_rsp_payload_transactionId, FetchPipelinePlugin_logic_retryIdCounter_value); // FetchPipelinePlugin2.scala:L448
              end
            `endif
          `endif
        end
      end
      if(FetchPipelinePlugin_logic_s4_logic_handleRsp) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((ICachePlugin_port_rsp_payload_transactionId == _zz_218)); // FetchPipelinePlugin2.scala:L454
          `else
            if(!(ICachePlugin_port_rsp_payload_transactionId == _zz_218)) begin
              $display("FAILURE ICache response TID mismatch! Expect %x, got %x", _zz_70, ICachePlugin_port_rsp_payload_transactionId); // FetchPipelinePlugin2.scala:L454
              $finish;
            end
          `endif
        `endif
        if(ICachePlugin_port_rsp_payload_redo) begin
          if(when_FetchPipelinePlugin2_l458) begin
            FetchPipelinePlugin_logic_retryCmd_lock <= 1'b1;
            FetchPipelinePlugin_logic_retryCmd_pc <= s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC;
            FetchPipelinePlugin_logic_retryCmd_id <= FetchPipelinePlugin_logic_retryIdCounter_value;
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // FetchPipelinePlugin2.scala:L464
              `else
                if(!1'b0) begin
                  $display("NOTE(FetchPipelinePlugin2.scala:464):  [notice] [33m[%x] FETCH-S4: Requesting retry for raw PC=0x%x, ID=%x, retryCmd.id=%x[0m", FetchPipelinePlugin_dbg_cycles, s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC, ICachePlugin_port_rsp_payload_transactionId, FetchPipelinePlugin_logic_retryIdCounter_value); // FetchPipelinePlugin2.scala:L464
                end
              `endif
            `endif
          end else begin
            if(when_FetchPipelinePlugin2_l467) begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // FetchPipelinePlugin2.scala:L468
                `else
                  if(!1'b0) begin
                    $display("NOTE(FetchPipelinePlugin2.scala:468):  [warning] [33m[%x] FETCH-S4: ICache requests retry for %x, but another retry for %x is already locked. Stalling.[0m", FetchPipelinePlugin_dbg_cycles, s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC, FetchPipelinePlugin_logic_retryCmd_pc); // FetchPipelinePlugin2.scala:L468
                  end
                `endif
              `endif
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // FetchPipelinePlugin2.scala:L469
                `else
                  if(!1'b0) begin
                    $display("FAILURE "); // FetchPipelinePlugin2.scala:L469
                    $finish;
                  end
                `endif
              `endif
            end
          end
        end else begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // FetchPipelinePlugin2.scala:L474
            `else
              if(!1'b0) begin
                $display("NOTE(FetchPipelinePlugin2.scala:474):  [success] [32m[%x] FETCH-S4: ICache hit for PC=0x%x[0m", FetchPipelinePlugin_dbg_cycles, s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC); // FetchPipelinePlugin2.scala:L474
              end
            `endif
          `endif
          if(when_FetchPipelinePlugin2_l476) begin
            FetchPipelinePlugin_logic_retryCmd_lock <= 1'b0;
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // FetchPipelinePlugin2.scala:L478
              `else
                if(!1'b0) begin
                  $display("NOTE(FetchPipelinePlugin2.scala:478):  [success] [32m[%x] FETCH-S4: Retry for ID %x completed. Clearing lock.[0m", FetchPipelinePlugin_dbg_cycles, FetchPipelinePlugin_logic_retryCmd_id); // FetchPipelinePlugin2.scala:L478
                end
              `endif
            `endif
          end
          if(when_FetchPipelinePlugin2_l481) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert((_zz_io_push_payload_numValidInstructions_1[1 : 0] == 2'b00)); // FetchPipelinePlugin2.scala:L166
              `else
                if(!(_zz_io_push_payload_numValidInstructions_1[1 : 0] == 2'b00)) begin
                  $display("FAILURE RAW_PC is not instruction-aligned within the cache line!"); // FetchPipelinePlugin2.scala:L166
                  $finish;
                end
              `endif
            `endif
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert((_zz_io_push_payload_numValidInstructions_1 < 32'h00000010)); // FetchPipelinePlugin2.scala:L168
              `else
                if(!(_zz_io_push_payload_numValidInstructions_1 < 32'h00000010)) begin
                  $display("FAILURE pcOffset exceeds cache line boundary!"); // FetchPipelinePlugin2.scala:L168
                  $finish;
                end
              `endif
            `endif
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(((! FetchPipelinePlugin_logic_doAnyFlush) && (! FetchPipelinePlugin_logic_isDrainingCacheRspReg))); // FetchPipelinePlugin2.scala:L501
              `else
                if(!((! FetchPipelinePlugin_logic_doAnyFlush) && (! FetchPipelinePlugin_logic_isDrainingCacheRspReg))) begin
                  $display("FAILURE Impossible to push valid predecoded group while flushing or draining cache Rsp."); // FetchPipelinePlugin2.scala:L501
                  $finish;
                end
              `endif
            `endif
            if(io_push_fire) begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // FetchPipelinePlugin2.scala:L507
                `else
                  if(!1'b0) begin
                    $display("NOTE(FetchPipelinePlugin2.scala:507):  [normal] FETCH-S4: Predecoded and pushing to FIFO. PC=0x%x, startIndex=%x, numValid=%x", s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC, _zz_io_push_payload_startInstructionIndex, _zz_io_push_payload_numValidInstructions); // FetchPipelinePlugin2.scala:L507
                  end
                `endif
              `endif
            end
          end
        end
      end
      if(io_fetchGroupIn_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L530
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:530):  [notice] [33m[DISPATCHER-IN] POP from predecodedGroups FIFO. PC=0x%x, startIdx=%x, numValid=%x, firstIsBranch=%x[0m", FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_pc, FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_startInstructionIndex, FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_pop_payload_numValidInstructions, _zz_71); // FetchPipelinePlugin2.scala:L530
            end
          `endif
        `endif
      end
      if(FetchPipelinePlugin_logic_s4_logic_predecodedGroups_io_flush) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L549
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:549):  [notice] [33m[%x] Flush predecodedGroups[0m", FetchPipelinePlugin_dbg_cycles); // FetchPipelinePlugin2.scala:L549
            end
          `endif
        `endif
      end
      if(FetchPipelinePlugin_logic_hardRedirect_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // FetchPipelinePlugin2.scala:L552
          `else
            if(!1'b0) begin
              $display("NOTE(FetchPipelinePlugin2.scala:552):  [notice] [33m[%x] Flush dispatcher[0m", FetchPipelinePlugin_dbg_cycles); // FetchPipelinePlugin2.scala:L552
            end
          `endif
        `endif
      end
      if(s1_PC_Gen_ready_output) begin
        s2_ICache_Access_valid <= _zz_s2_ICache_Access_valid;
      end
      if(when_Connection_l66_12) begin
        s2_ICache_Access_valid <= 1'b0;
      end
      if(s2_ICache_Access_ready_output) begin
        s4_Predecode_valid <= _zz_s4_Predecode_valid;
      end
      if(FetchPipelinePlugin_logic_hardRedirect_valid) begin
        s4_Predecode_valid <= 1'b0;
      end
      _zz_DataCachePlugin_logic_load_ohHistory_1 <= _zz_DataCachePlugin_logic_load_ohHistory_0;
      _zz_DataCachePlugin_logic_load_ohHistory_2 <= _zz_DataCachePlugin_logic_load_ohHistory_1;
      if(ROBPlugin_aggregatedFlushSignal_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // ROBPlugin.scala:L177
          `else
            if(!1'b0) begin
              $display("NOTE(ROBPlugin.scala:177):  [ROBPlugin] Aggregated flush signal is valid! Total ports: 1"); // ROBPlugin.scala:L177
            end
          `endif
        `endif
      end
      if(CommitPlugin_hw_robFlushPort_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // ROBPlugin.scala:L181
          `else
            if(!1'b0) begin
              $display("NOTE(ROBPlugin.scala:181):  [ROBPlugin] Flush port 0 is valid (reason=%s)", CommitPlugin_hw_robFlushPort_payload_reason_string); // ROBPlugin.scala:L181
            end
          `endif
        `endif
      end
      if(ROBPlugin_aggregatedFlushSignal_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // ROBPlugin.scala:L197
          `else
            if(!1'b0) begin
              $display("NOTE(ROBPlugin.scala:197):  [ROBPlugin] ROB component flush input is valid!"); // ROBPlugin.scala:L197
            end
          `endif
        `endif
      end
      if(when_CheckpointManagerPlugin_l117) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // CheckpointManagerPlugin.scala:L118
          `else
            if(!1'b0) begin
              $display("FAILURE Checkpoint restore requested but no valid checkpoint available"); // CheckpointManagerPlugin.scala:L118
              $finish;
            end
          `endif
        `endif
      end
      if(ICache_F1_Access_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_address[3 : 0] == 4'b0000)); // ICachePlugin.scala:L102
          `else
            if(!(ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_address[3 : 0] == 4'b0000)) begin
              $display("FAILURE ICache request must be line-aligned!"); // ICachePlugin.scala:L102
              $finish;
            end
          `endif
        `endif
      end
      ICachePlugin_logic_refill_refillCounter_value <= ICachePlugin_logic_refill_refillCounter_valueNext;
      ICachePlugin_logic_refill_fsm_stateReg <= ICachePlugin_logic_refill_fsm_stateNext;
      (* parallel_case *)
      case(1) // synthesis parallel_case
        (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
        end
        (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
        end
        (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
        end
        (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
          if(_zz_209[0]) begin
            if(_zz_81) begin
              ICachePlugin_logic_storage_valids_0_0 <= 1'b1;
            end
            if(_zz_82) begin
              ICachePlugin_logic_storage_valids_1_0 <= 1'b1;
            end
            if(_zz_83) begin
              ICachePlugin_logic_storage_valids_2_0 <= 1'b1;
            end
            if(_zz_84) begin
              ICachePlugin_logic_storage_valids_3_0 <= 1'b1;
            end
            if(_zz_85) begin
              ICachePlugin_logic_storage_valids_4_0 <= 1'b1;
            end
            if(_zz_86) begin
              ICachePlugin_logic_storage_valids_5_0 <= 1'b1;
            end
            if(_zz_87) begin
              ICachePlugin_logic_storage_valids_6_0 <= 1'b1;
            end
            if(_zz_88) begin
              ICachePlugin_logic_storage_valids_7_0 <= 1'b1;
            end
            if(_zz_89) begin
              ICachePlugin_logic_storage_valids_8_0 <= 1'b1;
            end
            if(_zz_90) begin
              ICachePlugin_logic_storage_valids_9_0 <= 1'b1;
            end
            if(_zz_91) begin
              ICachePlugin_logic_storage_valids_10_0 <= 1'b1;
            end
            if(_zz_92) begin
              ICachePlugin_logic_storage_valids_11_0 <= 1'b1;
            end
            if(_zz_93) begin
              ICachePlugin_logic_storage_valids_12_0 <= 1'b1;
            end
            if(_zz_94) begin
              ICachePlugin_logic_storage_valids_13_0 <= 1'b1;
            end
            if(_zz_95) begin
              ICachePlugin_logic_storage_valids_14_0 <= 1'b1;
            end
            if(_zz_96) begin
              ICachePlugin_logic_storage_valids_15_0 <= 1'b1;
            end
            if(_zz_97) begin
              ICachePlugin_logic_storage_valids_16_0 <= 1'b1;
            end
            if(_zz_98) begin
              ICachePlugin_logic_storage_valids_17_0 <= 1'b1;
            end
            if(_zz_99) begin
              ICachePlugin_logic_storage_valids_18_0 <= 1'b1;
            end
            if(_zz_100) begin
              ICachePlugin_logic_storage_valids_19_0 <= 1'b1;
            end
            if(_zz_101) begin
              ICachePlugin_logic_storage_valids_20_0 <= 1'b1;
            end
            if(_zz_102) begin
              ICachePlugin_logic_storage_valids_21_0 <= 1'b1;
            end
            if(_zz_103) begin
              ICachePlugin_logic_storage_valids_22_0 <= 1'b1;
            end
            if(_zz_104) begin
              ICachePlugin_logic_storage_valids_23_0 <= 1'b1;
            end
            if(_zz_105) begin
              ICachePlugin_logic_storage_valids_24_0 <= 1'b1;
            end
            if(_zz_106) begin
              ICachePlugin_logic_storage_valids_25_0 <= 1'b1;
            end
            if(_zz_107) begin
              ICachePlugin_logic_storage_valids_26_0 <= 1'b1;
            end
            if(_zz_108) begin
              ICachePlugin_logic_storage_valids_27_0 <= 1'b1;
            end
            if(_zz_109) begin
              ICachePlugin_logic_storage_valids_28_0 <= 1'b1;
            end
            if(_zz_110) begin
              ICachePlugin_logic_storage_valids_29_0 <= 1'b1;
            end
            if(_zz_111) begin
              ICachePlugin_logic_storage_valids_30_0 <= 1'b1;
            end
            if(_zz_112) begin
              ICachePlugin_logic_storage_valids_31_0 <= 1'b1;
            end
            if(_zz_113) begin
              ICachePlugin_logic_storage_valids_32_0 <= 1'b1;
            end
            if(_zz_114) begin
              ICachePlugin_logic_storage_valids_33_0 <= 1'b1;
            end
            if(_zz_115) begin
              ICachePlugin_logic_storage_valids_34_0 <= 1'b1;
            end
            if(_zz_116) begin
              ICachePlugin_logic_storage_valids_35_0 <= 1'b1;
            end
            if(_zz_117) begin
              ICachePlugin_logic_storage_valids_36_0 <= 1'b1;
            end
            if(_zz_118) begin
              ICachePlugin_logic_storage_valids_37_0 <= 1'b1;
            end
            if(_zz_119) begin
              ICachePlugin_logic_storage_valids_38_0 <= 1'b1;
            end
            if(_zz_120) begin
              ICachePlugin_logic_storage_valids_39_0 <= 1'b1;
            end
            if(_zz_121) begin
              ICachePlugin_logic_storage_valids_40_0 <= 1'b1;
            end
            if(_zz_122) begin
              ICachePlugin_logic_storage_valids_41_0 <= 1'b1;
            end
            if(_zz_123) begin
              ICachePlugin_logic_storage_valids_42_0 <= 1'b1;
            end
            if(_zz_124) begin
              ICachePlugin_logic_storage_valids_43_0 <= 1'b1;
            end
            if(_zz_125) begin
              ICachePlugin_logic_storage_valids_44_0 <= 1'b1;
            end
            if(_zz_126) begin
              ICachePlugin_logic_storage_valids_45_0 <= 1'b1;
            end
            if(_zz_127) begin
              ICachePlugin_logic_storage_valids_46_0 <= 1'b1;
            end
            if(_zz_128) begin
              ICachePlugin_logic_storage_valids_47_0 <= 1'b1;
            end
            if(_zz_129) begin
              ICachePlugin_logic_storage_valids_48_0 <= 1'b1;
            end
            if(_zz_130) begin
              ICachePlugin_logic_storage_valids_49_0 <= 1'b1;
            end
            if(_zz_131) begin
              ICachePlugin_logic_storage_valids_50_0 <= 1'b1;
            end
            if(_zz_132) begin
              ICachePlugin_logic_storage_valids_51_0 <= 1'b1;
            end
            if(_zz_133) begin
              ICachePlugin_logic_storage_valids_52_0 <= 1'b1;
            end
            if(_zz_134) begin
              ICachePlugin_logic_storage_valids_53_0 <= 1'b1;
            end
            if(_zz_135) begin
              ICachePlugin_logic_storage_valids_54_0 <= 1'b1;
            end
            if(_zz_136) begin
              ICachePlugin_logic_storage_valids_55_0 <= 1'b1;
            end
            if(_zz_137) begin
              ICachePlugin_logic_storage_valids_56_0 <= 1'b1;
            end
            if(_zz_138) begin
              ICachePlugin_logic_storage_valids_57_0 <= 1'b1;
            end
            if(_zz_139) begin
              ICachePlugin_logic_storage_valids_58_0 <= 1'b1;
            end
            if(_zz_140) begin
              ICachePlugin_logic_storage_valids_59_0 <= 1'b1;
            end
            if(_zz_141) begin
              ICachePlugin_logic_storage_valids_60_0 <= 1'b1;
            end
            if(_zz_142) begin
              ICachePlugin_logic_storage_valids_61_0 <= 1'b1;
            end
            if(_zz_143) begin
              ICachePlugin_logic_storage_valids_62_0 <= 1'b1;
            end
            if(_zz_144) begin
              ICachePlugin_logic_storage_valids_63_0 <= 1'b1;
            end
            if(_zz_145) begin
              ICachePlugin_logic_storage_valids_64_0 <= 1'b1;
            end
            if(_zz_146) begin
              ICachePlugin_logic_storage_valids_65_0 <= 1'b1;
            end
            if(_zz_147) begin
              ICachePlugin_logic_storage_valids_66_0 <= 1'b1;
            end
            if(_zz_148) begin
              ICachePlugin_logic_storage_valids_67_0 <= 1'b1;
            end
            if(_zz_149) begin
              ICachePlugin_logic_storage_valids_68_0 <= 1'b1;
            end
            if(_zz_150) begin
              ICachePlugin_logic_storage_valids_69_0 <= 1'b1;
            end
            if(_zz_151) begin
              ICachePlugin_logic_storage_valids_70_0 <= 1'b1;
            end
            if(_zz_152) begin
              ICachePlugin_logic_storage_valids_71_0 <= 1'b1;
            end
            if(_zz_153) begin
              ICachePlugin_logic_storage_valids_72_0 <= 1'b1;
            end
            if(_zz_154) begin
              ICachePlugin_logic_storage_valids_73_0 <= 1'b1;
            end
            if(_zz_155) begin
              ICachePlugin_logic_storage_valids_74_0 <= 1'b1;
            end
            if(_zz_156) begin
              ICachePlugin_logic_storage_valids_75_0 <= 1'b1;
            end
            if(_zz_157) begin
              ICachePlugin_logic_storage_valids_76_0 <= 1'b1;
            end
            if(_zz_158) begin
              ICachePlugin_logic_storage_valids_77_0 <= 1'b1;
            end
            if(_zz_159) begin
              ICachePlugin_logic_storage_valids_78_0 <= 1'b1;
            end
            if(_zz_160) begin
              ICachePlugin_logic_storage_valids_79_0 <= 1'b1;
            end
            if(_zz_161) begin
              ICachePlugin_logic_storage_valids_80_0 <= 1'b1;
            end
            if(_zz_162) begin
              ICachePlugin_logic_storage_valids_81_0 <= 1'b1;
            end
            if(_zz_163) begin
              ICachePlugin_logic_storage_valids_82_0 <= 1'b1;
            end
            if(_zz_164) begin
              ICachePlugin_logic_storage_valids_83_0 <= 1'b1;
            end
            if(_zz_165) begin
              ICachePlugin_logic_storage_valids_84_0 <= 1'b1;
            end
            if(_zz_166) begin
              ICachePlugin_logic_storage_valids_85_0 <= 1'b1;
            end
            if(_zz_167) begin
              ICachePlugin_logic_storage_valids_86_0 <= 1'b1;
            end
            if(_zz_168) begin
              ICachePlugin_logic_storage_valids_87_0 <= 1'b1;
            end
            if(_zz_169) begin
              ICachePlugin_logic_storage_valids_88_0 <= 1'b1;
            end
            if(_zz_170) begin
              ICachePlugin_logic_storage_valids_89_0 <= 1'b1;
            end
            if(_zz_171) begin
              ICachePlugin_logic_storage_valids_90_0 <= 1'b1;
            end
            if(_zz_172) begin
              ICachePlugin_logic_storage_valids_91_0 <= 1'b1;
            end
            if(_zz_173) begin
              ICachePlugin_logic_storage_valids_92_0 <= 1'b1;
            end
            if(_zz_174) begin
              ICachePlugin_logic_storage_valids_93_0 <= 1'b1;
            end
            if(_zz_175) begin
              ICachePlugin_logic_storage_valids_94_0 <= 1'b1;
            end
            if(_zz_176) begin
              ICachePlugin_logic_storage_valids_95_0 <= 1'b1;
            end
            if(_zz_177) begin
              ICachePlugin_logic_storage_valids_96_0 <= 1'b1;
            end
            if(_zz_178) begin
              ICachePlugin_logic_storage_valids_97_0 <= 1'b1;
            end
            if(_zz_179) begin
              ICachePlugin_logic_storage_valids_98_0 <= 1'b1;
            end
            if(_zz_180) begin
              ICachePlugin_logic_storage_valids_99_0 <= 1'b1;
            end
            if(_zz_181) begin
              ICachePlugin_logic_storage_valids_100_0 <= 1'b1;
            end
            if(_zz_182) begin
              ICachePlugin_logic_storage_valids_101_0 <= 1'b1;
            end
            if(_zz_183) begin
              ICachePlugin_logic_storage_valids_102_0 <= 1'b1;
            end
            if(_zz_184) begin
              ICachePlugin_logic_storage_valids_103_0 <= 1'b1;
            end
            if(_zz_185) begin
              ICachePlugin_logic_storage_valids_104_0 <= 1'b1;
            end
            if(_zz_186) begin
              ICachePlugin_logic_storage_valids_105_0 <= 1'b1;
            end
            if(_zz_187) begin
              ICachePlugin_logic_storage_valids_106_0 <= 1'b1;
            end
            if(_zz_188) begin
              ICachePlugin_logic_storage_valids_107_0 <= 1'b1;
            end
            if(_zz_189) begin
              ICachePlugin_logic_storage_valids_108_0 <= 1'b1;
            end
            if(_zz_190) begin
              ICachePlugin_logic_storage_valids_109_0 <= 1'b1;
            end
            if(_zz_191) begin
              ICachePlugin_logic_storage_valids_110_0 <= 1'b1;
            end
            if(_zz_192) begin
              ICachePlugin_logic_storage_valids_111_0 <= 1'b1;
            end
            if(_zz_193) begin
              ICachePlugin_logic_storage_valids_112_0 <= 1'b1;
            end
            if(_zz_194) begin
              ICachePlugin_logic_storage_valids_113_0 <= 1'b1;
            end
            if(_zz_195) begin
              ICachePlugin_logic_storage_valids_114_0 <= 1'b1;
            end
            if(_zz_196) begin
              ICachePlugin_logic_storage_valids_115_0 <= 1'b1;
            end
            if(_zz_197) begin
              ICachePlugin_logic_storage_valids_116_0 <= 1'b1;
            end
            if(_zz_198) begin
              ICachePlugin_logic_storage_valids_117_0 <= 1'b1;
            end
            if(_zz_199) begin
              ICachePlugin_logic_storage_valids_118_0 <= 1'b1;
            end
            if(_zz_200) begin
              ICachePlugin_logic_storage_valids_119_0 <= 1'b1;
            end
            if(_zz_201) begin
              ICachePlugin_logic_storage_valids_120_0 <= 1'b1;
            end
            if(_zz_202) begin
              ICachePlugin_logic_storage_valids_121_0 <= 1'b1;
            end
            if(_zz_203) begin
              ICachePlugin_logic_storage_valids_122_0 <= 1'b1;
            end
            if(_zz_204) begin
              ICachePlugin_logic_storage_valids_123_0 <= 1'b1;
            end
            if(_zz_205) begin
              ICachePlugin_logic_storage_valids_124_0 <= 1'b1;
            end
            if(_zz_206) begin
              ICachePlugin_logic_storage_valids_125_0 <= 1'b1;
            end
            if(_zz_207) begin
              ICachePlugin_logic_storage_valids_126_0 <= 1'b1;
            end
            if(_zz_208) begin
              ICachePlugin_logic_storage_valids_127_0 <= 1'b1;
            end
          end
          if(_zz_209[1]) begin
            if(_zz_81) begin
              ICachePlugin_logic_storage_valids_0_1 <= 1'b1;
            end
            if(_zz_82) begin
              ICachePlugin_logic_storage_valids_1_1 <= 1'b1;
            end
            if(_zz_83) begin
              ICachePlugin_logic_storage_valids_2_1 <= 1'b1;
            end
            if(_zz_84) begin
              ICachePlugin_logic_storage_valids_3_1 <= 1'b1;
            end
            if(_zz_85) begin
              ICachePlugin_logic_storage_valids_4_1 <= 1'b1;
            end
            if(_zz_86) begin
              ICachePlugin_logic_storage_valids_5_1 <= 1'b1;
            end
            if(_zz_87) begin
              ICachePlugin_logic_storage_valids_6_1 <= 1'b1;
            end
            if(_zz_88) begin
              ICachePlugin_logic_storage_valids_7_1 <= 1'b1;
            end
            if(_zz_89) begin
              ICachePlugin_logic_storage_valids_8_1 <= 1'b1;
            end
            if(_zz_90) begin
              ICachePlugin_logic_storage_valids_9_1 <= 1'b1;
            end
            if(_zz_91) begin
              ICachePlugin_logic_storage_valids_10_1 <= 1'b1;
            end
            if(_zz_92) begin
              ICachePlugin_logic_storage_valids_11_1 <= 1'b1;
            end
            if(_zz_93) begin
              ICachePlugin_logic_storage_valids_12_1 <= 1'b1;
            end
            if(_zz_94) begin
              ICachePlugin_logic_storage_valids_13_1 <= 1'b1;
            end
            if(_zz_95) begin
              ICachePlugin_logic_storage_valids_14_1 <= 1'b1;
            end
            if(_zz_96) begin
              ICachePlugin_logic_storage_valids_15_1 <= 1'b1;
            end
            if(_zz_97) begin
              ICachePlugin_logic_storage_valids_16_1 <= 1'b1;
            end
            if(_zz_98) begin
              ICachePlugin_logic_storage_valids_17_1 <= 1'b1;
            end
            if(_zz_99) begin
              ICachePlugin_logic_storage_valids_18_1 <= 1'b1;
            end
            if(_zz_100) begin
              ICachePlugin_logic_storage_valids_19_1 <= 1'b1;
            end
            if(_zz_101) begin
              ICachePlugin_logic_storage_valids_20_1 <= 1'b1;
            end
            if(_zz_102) begin
              ICachePlugin_logic_storage_valids_21_1 <= 1'b1;
            end
            if(_zz_103) begin
              ICachePlugin_logic_storage_valids_22_1 <= 1'b1;
            end
            if(_zz_104) begin
              ICachePlugin_logic_storage_valids_23_1 <= 1'b1;
            end
            if(_zz_105) begin
              ICachePlugin_logic_storage_valids_24_1 <= 1'b1;
            end
            if(_zz_106) begin
              ICachePlugin_logic_storage_valids_25_1 <= 1'b1;
            end
            if(_zz_107) begin
              ICachePlugin_logic_storage_valids_26_1 <= 1'b1;
            end
            if(_zz_108) begin
              ICachePlugin_logic_storage_valids_27_1 <= 1'b1;
            end
            if(_zz_109) begin
              ICachePlugin_logic_storage_valids_28_1 <= 1'b1;
            end
            if(_zz_110) begin
              ICachePlugin_logic_storage_valids_29_1 <= 1'b1;
            end
            if(_zz_111) begin
              ICachePlugin_logic_storage_valids_30_1 <= 1'b1;
            end
            if(_zz_112) begin
              ICachePlugin_logic_storage_valids_31_1 <= 1'b1;
            end
            if(_zz_113) begin
              ICachePlugin_logic_storage_valids_32_1 <= 1'b1;
            end
            if(_zz_114) begin
              ICachePlugin_logic_storage_valids_33_1 <= 1'b1;
            end
            if(_zz_115) begin
              ICachePlugin_logic_storage_valids_34_1 <= 1'b1;
            end
            if(_zz_116) begin
              ICachePlugin_logic_storage_valids_35_1 <= 1'b1;
            end
            if(_zz_117) begin
              ICachePlugin_logic_storage_valids_36_1 <= 1'b1;
            end
            if(_zz_118) begin
              ICachePlugin_logic_storage_valids_37_1 <= 1'b1;
            end
            if(_zz_119) begin
              ICachePlugin_logic_storage_valids_38_1 <= 1'b1;
            end
            if(_zz_120) begin
              ICachePlugin_logic_storage_valids_39_1 <= 1'b1;
            end
            if(_zz_121) begin
              ICachePlugin_logic_storage_valids_40_1 <= 1'b1;
            end
            if(_zz_122) begin
              ICachePlugin_logic_storage_valids_41_1 <= 1'b1;
            end
            if(_zz_123) begin
              ICachePlugin_logic_storage_valids_42_1 <= 1'b1;
            end
            if(_zz_124) begin
              ICachePlugin_logic_storage_valids_43_1 <= 1'b1;
            end
            if(_zz_125) begin
              ICachePlugin_logic_storage_valids_44_1 <= 1'b1;
            end
            if(_zz_126) begin
              ICachePlugin_logic_storage_valids_45_1 <= 1'b1;
            end
            if(_zz_127) begin
              ICachePlugin_logic_storage_valids_46_1 <= 1'b1;
            end
            if(_zz_128) begin
              ICachePlugin_logic_storage_valids_47_1 <= 1'b1;
            end
            if(_zz_129) begin
              ICachePlugin_logic_storage_valids_48_1 <= 1'b1;
            end
            if(_zz_130) begin
              ICachePlugin_logic_storage_valids_49_1 <= 1'b1;
            end
            if(_zz_131) begin
              ICachePlugin_logic_storage_valids_50_1 <= 1'b1;
            end
            if(_zz_132) begin
              ICachePlugin_logic_storage_valids_51_1 <= 1'b1;
            end
            if(_zz_133) begin
              ICachePlugin_logic_storage_valids_52_1 <= 1'b1;
            end
            if(_zz_134) begin
              ICachePlugin_logic_storage_valids_53_1 <= 1'b1;
            end
            if(_zz_135) begin
              ICachePlugin_logic_storage_valids_54_1 <= 1'b1;
            end
            if(_zz_136) begin
              ICachePlugin_logic_storage_valids_55_1 <= 1'b1;
            end
            if(_zz_137) begin
              ICachePlugin_logic_storage_valids_56_1 <= 1'b1;
            end
            if(_zz_138) begin
              ICachePlugin_logic_storage_valids_57_1 <= 1'b1;
            end
            if(_zz_139) begin
              ICachePlugin_logic_storage_valids_58_1 <= 1'b1;
            end
            if(_zz_140) begin
              ICachePlugin_logic_storage_valids_59_1 <= 1'b1;
            end
            if(_zz_141) begin
              ICachePlugin_logic_storage_valids_60_1 <= 1'b1;
            end
            if(_zz_142) begin
              ICachePlugin_logic_storage_valids_61_1 <= 1'b1;
            end
            if(_zz_143) begin
              ICachePlugin_logic_storage_valids_62_1 <= 1'b1;
            end
            if(_zz_144) begin
              ICachePlugin_logic_storage_valids_63_1 <= 1'b1;
            end
            if(_zz_145) begin
              ICachePlugin_logic_storage_valids_64_1 <= 1'b1;
            end
            if(_zz_146) begin
              ICachePlugin_logic_storage_valids_65_1 <= 1'b1;
            end
            if(_zz_147) begin
              ICachePlugin_logic_storage_valids_66_1 <= 1'b1;
            end
            if(_zz_148) begin
              ICachePlugin_logic_storage_valids_67_1 <= 1'b1;
            end
            if(_zz_149) begin
              ICachePlugin_logic_storage_valids_68_1 <= 1'b1;
            end
            if(_zz_150) begin
              ICachePlugin_logic_storage_valids_69_1 <= 1'b1;
            end
            if(_zz_151) begin
              ICachePlugin_logic_storage_valids_70_1 <= 1'b1;
            end
            if(_zz_152) begin
              ICachePlugin_logic_storage_valids_71_1 <= 1'b1;
            end
            if(_zz_153) begin
              ICachePlugin_logic_storage_valids_72_1 <= 1'b1;
            end
            if(_zz_154) begin
              ICachePlugin_logic_storage_valids_73_1 <= 1'b1;
            end
            if(_zz_155) begin
              ICachePlugin_logic_storage_valids_74_1 <= 1'b1;
            end
            if(_zz_156) begin
              ICachePlugin_logic_storage_valids_75_1 <= 1'b1;
            end
            if(_zz_157) begin
              ICachePlugin_logic_storage_valids_76_1 <= 1'b1;
            end
            if(_zz_158) begin
              ICachePlugin_logic_storage_valids_77_1 <= 1'b1;
            end
            if(_zz_159) begin
              ICachePlugin_logic_storage_valids_78_1 <= 1'b1;
            end
            if(_zz_160) begin
              ICachePlugin_logic_storage_valids_79_1 <= 1'b1;
            end
            if(_zz_161) begin
              ICachePlugin_logic_storage_valids_80_1 <= 1'b1;
            end
            if(_zz_162) begin
              ICachePlugin_logic_storage_valids_81_1 <= 1'b1;
            end
            if(_zz_163) begin
              ICachePlugin_logic_storage_valids_82_1 <= 1'b1;
            end
            if(_zz_164) begin
              ICachePlugin_logic_storage_valids_83_1 <= 1'b1;
            end
            if(_zz_165) begin
              ICachePlugin_logic_storage_valids_84_1 <= 1'b1;
            end
            if(_zz_166) begin
              ICachePlugin_logic_storage_valids_85_1 <= 1'b1;
            end
            if(_zz_167) begin
              ICachePlugin_logic_storage_valids_86_1 <= 1'b1;
            end
            if(_zz_168) begin
              ICachePlugin_logic_storage_valids_87_1 <= 1'b1;
            end
            if(_zz_169) begin
              ICachePlugin_logic_storage_valids_88_1 <= 1'b1;
            end
            if(_zz_170) begin
              ICachePlugin_logic_storage_valids_89_1 <= 1'b1;
            end
            if(_zz_171) begin
              ICachePlugin_logic_storage_valids_90_1 <= 1'b1;
            end
            if(_zz_172) begin
              ICachePlugin_logic_storage_valids_91_1 <= 1'b1;
            end
            if(_zz_173) begin
              ICachePlugin_logic_storage_valids_92_1 <= 1'b1;
            end
            if(_zz_174) begin
              ICachePlugin_logic_storage_valids_93_1 <= 1'b1;
            end
            if(_zz_175) begin
              ICachePlugin_logic_storage_valids_94_1 <= 1'b1;
            end
            if(_zz_176) begin
              ICachePlugin_logic_storage_valids_95_1 <= 1'b1;
            end
            if(_zz_177) begin
              ICachePlugin_logic_storage_valids_96_1 <= 1'b1;
            end
            if(_zz_178) begin
              ICachePlugin_logic_storage_valids_97_1 <= 1'b1;
            end
            if(_zz_179) begin
              ICachePlugin_logic_storage_valids_98_1 <= 1'b1;
            end
            if(_zz_180) begin
              ICachePlugin_logic_storage_valids_99_1 <= 1'b1;
            end
            if(_zz_181) begin
              ICachePlugin_logic_storage_valids_100_1 <= 1'b1;
            end
            if(_zz_182) begin
              ICachePlugin_logic_storage_valids_101_1 <= 1'b1;
            end
            if(_zz_183) begin
              ICachePlugin_logic_storage_valids_102_1 <= 1'b1;
            end
            if(_zz_184) begin
              ICachePlugin_logic_storage_valids_103_1 <= 1'b1;
            end
            if(_zz_185) begin
              ICachePlugin_logic_storage_valids_104_1 <= 1'b1;
            end
            if(_zz_186) begin
              ICachePlugin_logic_storage_valids_105_1 <= 1'b1;
            end
            if(_zz_187) begin
              ICachePlugin_logic_storage_valids_106_1 <= 1'b1;
            end
            if(_zz_188) begin
              ICachePlugin_logic_storage_valids_107_1 <= 1'b1;
            end
            if(_zz_189) begin
              ICachePlugin_logic_storage_valids_108_1 <= 1'b1;
            end
            if(_zz_190) begin
              ICachePlugin_logic_storage_valids_109_1 <= 1'b1;
            end
            if(_zz_191) begin
              ICachePlugin_logic_storage_valids_110_1 <= 1'b1;
            end
            if(_zz_192) begin
              ICachePlugin_logic_storage_valids_111_1 <= 1'b1;
            end
            if(_zz_193) begin
              ICachePlugin_logic_storage_valids_112_1 <= 1'b1;
            end
            if(_zz_194) begin
              ICachePlugin_logic_storage_valids_113_1 <= 1'b1;
            end
            if(_zz_195) begin
              ICachePlugin_logic_storage_valids_114_1 <= 1'b1;
            end
            if(_zz_196) begin
              ICachePlugin_logic_storage_valids_115_1 <= 1'b1;
            end
            if(_zz_197) begin
              ICachePlugin_logic_storage_valids_116_1 <= 1'b1;
            end
            if(_zz_198) begin
              ICachePlugin_logic_storage_valids_117_1 <= 1'b1;
            end
            if(_zz_199) begin
              ICachePlugin_logic_storage_valids_118_1 <= 1'b1;
            end
            if(_zz_200) begin
              ICachePlugin_logic_storage_valids_119_1 <= 1'b1;
            end
            if(_zz_201) begin
              ICachePlugin_logic_storage_valids_120_1 <= 1'b1;
            end
            if(_zz_202) begin
              ICachePlugin_logic_storage_valids_121_1 <= 1'b1;
            end
            if(_zz_203) begin
              ICachePlugin_logic_storage_valids_122_1 <= 1'b1;
            end
            if(_zz_204) begin
              ICachePlugin_logic_storage_valids_123_1 <= 1'b1;
            end
            if(_zz_205) begin
              ICachePlugin_logic_storage_valids_124_1 <= 1'b1;
            end
            if(_zz_206) begin
              ICachePlugin_logic_storage_valids_125_1 <= 1'b1;
            end
            if(_zz_207) begin
              ICachePlugin_logic_storage_valids_126_1 <= 1'b1;
            end
            if(_zz_208) begin
              ICachePlugin_logic_storage_valids_127_1 <= 1'b1;
            end
          end
        end
        default : begin
        end
      endcase
      if(ICachePlugin_invalidate) begin
        ICachePlugin_logic_storage_valids_0_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_0_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_1_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_1_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_2_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_2_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_3_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_3_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_4_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_4_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_5_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_5_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_6_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_6_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_7_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_7_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_8_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_8_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_9_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_9_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_10_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_10_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_11_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_11_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_12_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_12_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_13_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_13_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_14_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_14_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_15_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_15_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_16_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_16_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_17_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_17_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_18_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_18_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_19_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_19_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_20_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_20_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_21_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_21_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_22_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_22_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_23_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_23_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_24_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_24_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_25_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_25_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_26_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_26_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_27_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_27_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_28_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_28_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_29_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_29_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_30_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_30_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_31_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_31_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_32_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_32_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_33_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_33_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_34_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_34_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_35_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_35_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_36_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_36_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_37_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_37_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_38_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_38_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_39_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_39_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_40_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_40_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_41_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_41_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_42_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_42_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_43_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_43_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_44_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_44_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_45_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_45_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_46_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_46_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_47_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_47_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_48_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_48_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_49_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_49_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_50_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_50_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_51_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_51_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_52_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_52_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_53_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_53_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_54_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_54_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_55_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_55_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_56_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_56_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_57_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_57_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_58_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_58_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_59_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_59_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_60_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_60_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_61_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_61_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_62_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_62_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_63_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_63_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_64_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_64_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_65_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_65_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_66_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_66_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_67_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_67_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_68_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_68_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_69_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_69_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_70_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_70_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_71_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_71_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_72_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_72_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_73_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_73_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_74_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_74_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_75_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_75_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_76_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_76_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_77_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_77_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_78_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_78_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_79_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_79_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_80_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_80_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_81_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_81_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_82_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_82_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_83_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_83_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_84_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_84_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_85_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_85_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_86_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_86_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_87_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_87_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_88_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_88_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_89_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_89_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_90_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_90_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_91_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_91_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_92_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_92_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_93_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_93_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_94_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_94_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_95_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_95_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_96_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_96_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_97_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_97_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_98_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_98_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_99_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_99_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_100_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_100_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_101_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_101_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_102_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_102_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_103_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_103_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_104_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_104_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_105_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_105_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_106_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_106_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_107_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_107_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_108_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_108_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_109_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_109_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_110_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_110_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_111_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_111_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_112_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_112_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_113_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_113_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_114_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_114_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_115_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_115_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_116_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_116_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_117_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_117_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_118_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_118_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_119_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_119_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_120_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_120_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_121_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_121_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_122_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_122_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_123_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_123_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_124_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_124_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_125_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_125_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_126_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_126_1 <= 1'b0;
        ICachePlugin_logic_storage_valids_127_0 <= 1'b0;
        ICachePlugin_logic_storage_valids_127_1 <= 1'b0;
      end
      ICache_F2_HitCheck_valid <= ICache_F1_Access_valid;
      if(BpuPipelinePlugin_logic_s1_read_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BpuPlugin.scala:L85
          `else
            if(!1'b0) begin
              $display("NOTE(BpuPlugin.scala:85):  [debug] [34m[BPU.S1] Query Firing for PC=0x%x, TID=%x, PHT Idx=0x%x, BTB Idx=0x%x[0m", BpuPipelinePlugin_logic_s1_read_Q_PC, BpuPipelinePlugin_logic_s1_read_TRANSACTION_ID, _zz_210, _zz_211); // BpuPlugin.scala:L85
            end
          `endif
        `endif
      end
      if(BpuPipelinePlugin_logic_s2_predict_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BpuPlugin.scala:L107
          `else
            if(!1'b0) begin
              $display("NOTE(BpuPlugin.scala:107):  [debug] [34m[BPU.S2] Predict Firing for PC=0x%x, TID=%x | PHT Readout=%x -> Predict=%x | BTB Readout: valid=%x tag_match=%x -> Hit=%x | Final Predict: isTaken=%x target=0x%x[0m", BpuPipelinePlugin_logic_s2_predict_Q_PC, BpuPipelinePlugin_logic_s2_predict_TRANSACTION_ID, BpuPipelinePlugin_logic_phtReadData_s1, BpuPipelinePlugin_logic_phtPrediction, BpuPipelinePlugin_logic_btbReadData_s1_valid, _zz_214, BpuPipelinePlugin_logic_btbHit, BpuPipelinePlugin_logic_s2_predict_IS_TAKEN, BpuPipelinePlugin_logic_s2_predict_TARGET_PC); // BpuPlugin.scala:L107
            end
          `endif
        `endif
      end
      if(BpuPipelinePlugin_logic_u1_read_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BpuPlugin.scala:L131
          `else
            if(!1'b0) begin
              $display("NOTE(BpuPlugin.scala:131):  [debug] [34m[BPU.U1] Update Firing for PC=0x%x, isTaken=%x[0m", BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_pc, BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_isTaken); // BpuPlugin.scala:L131
            end
          `endif
        `endif
      end
      if(BpuPipelinePlugin_logic_u2_write_isFiring) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BpuPlugin.scala:L152
          `else
            if(!1'b0) begin
              $display("NOTE(BpuPlugin.scala:152):  [debug] [34m[BPU.U2] Write Firing for PC=0x%x | Old PHT=%x -> New PHT=%x | isTaken=%x, Wr BTB?=%x[0m", BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_pc, BpuPipelinePlugin_logic_oldPhtState_u1, BpuPipelinePlugin_logic_newPhtState, BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken, BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken); // BpuPlugin.scala:L152
            end
          `endif
        `endif
      end
      if(BpuPipelinePlugin_logic_s2_predict_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BpuPlugin.scala:L230
          `else
            if(!1'b0) begin
              $display("NOTE(BpuPlugin.scala:230):  [BPU] Query PC=0x%x, TID=%x -> Predict: isTaken=%x target=0x%x", BpuPipelinePlugin_queryPortIn_payload_pc_regNext, BpuPipelinePlugin_queryPortIn_payload_transactionId_regNext, BpuPipelinePlugin_responseFlowOut_payload_isTaken, BpuPipelinePlugin_responseFlowOut_payload_target); // BpuPlugin.scala:L230
            end
          `endif
        `endif
      end
      BpuPipelinePlugin_logic_s2_predict_valid <= BpuPipelinePlugin_logic_s1_read_valid;
      BpuPipelinePlugin_logic_u2_write_valid <= BpuPipelinePlugin_logic_u1_read_valid;
      if(FetchPipelinePlugin_doHardRedirect_listening) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // BpuPlugin.scala:L251
          `else
            if(!1'b0) begin
              $display("NOTE(BpuPlugin.scala:251):  [BPU] FLUSH: Flushing internal query and update pipelines due to hard redirect."); // BpuPlugin.scala:L251
            end
          `endif
        `endif
      end
      if(io_axiOut_readOnly_decoder_io_outputs_0_ar_valid) begin
        io_outputs_0_ar_rValid <= 1'b1;
      end
      if(io_outputs_0_ar_validPipe_fire) begin
        io_outputs_0_ar_rValid <= 1'b0;
      end
      if(io_axiOut_readOnly_decoder_io_outputs_1_ar_valid) begin
        io_outputs_1_ar_rValid <= 1'b1;
      end
      if(io_outputs_1_ar_validPipe_fire) begin
        io_outputs_1_ar_rValid <= 1'b0;
      end
      if(io_axiOut_readOnly_decoder_io_outputs_2_ar_valid) begin
        io_outputs_2_ar_rValid <= 1'b1;
      end
      if(io_outputs_2_ar_validPipe_fire) begin
        io_outputs_2_ar_rValid <= 1'b0;
      end
      if(io_axiOut_writeOnly_decoder_io_outputs_0_aw_valid) begin
        io_outputs_0_aw_rValid <= 1'b1;
      end
      if(io_outputs_0_aw_validPipe_fire) begin
        io_outputs_0_aw_rValid <= 1'b0;
      end
      if(io_axiOut_writeOnly_decoder_io_outputs_1_aw_valid) begin
        io_outputs_1_aw_rValid <= 1'b1;
      end
      if(io_outputs_1_aw_validPipe_fire) begin
        io_outputs_1_aw_rValid <= 1'b0;
      end
      if(io_axiOut_writeOnly_decoder_io_outputs_2_aw_valid) begin
        io_outputs_2_aw_rValid <= 1'b1;
      end
      if(io_outputs_2_aw_validPipe_fire) begin
        io_outputs_2_aw_rValid <= 1'b0;
      end
      if(io_axiOut_readOnly_decoder_1_io_outputs_0_ar_valid) begin
        io_outputs_0_ar_rValid_1 <= 1'b1;
      end
      if(io_outputs_0_ar_validPipe_fire_1) begin
        io_outputs_0_ar_rValid_1 <= 1'b0;
      end
      if(io_axiOut_readOnly_decoder_1_io_outputs_1_ar_valid) begin
        io_outputs_1_ar_rValid_1 <= 1'b1;
      end
      if(io_outputs_1_ar_validPipe_fire_1) begin
        io_outputs_1_ar_rValid_1 <= 1'b0;
      end
      if(io_axiOut_readOnly_decoder_1_io_outputs_2_ar_valid) begin
        io_outputs_2_ar_rValid_1 <= 1'b1;
      end
      if(io_outputs_2_ar_validPipe_fire_1) begin
        io_outputs_2_ar_rValid_1 <= 1'b0;
      end
      if(io_axiOut_writeOnly_decoder_1_io_outputs_0_aw_valid) begin
        io_outputs_0_aw_rValid_1 <= 1'b1;
      end
      if(io_outputs_0_aw_validPipe_fire_1) begin
        io_outputs_0_aw_rValid_1 <= 1'b0;
      end
      if(io_axiOut_writeOnly_decoder_1_io_outputs_1_aw_valid) begin
        io_outputs_1_aw_rValid_1 <= 1'b1;
      end
      if(io_outputs_1_aw_validPipe_fire_1) begin
        io_outputs_1_aw_rValid_1 <= 1'b0;
      end
      if(io_axiOut_writeOnly_decoder_1_io_outputs_2_aw_valid) begin
        io_outputs_2_aw_rValid_1 <= 1'b1;
      end
      if(io_outputs_2_aw_validPipe_fire_1) begin
        io_outputs_2_aw_rValid_1 <= 1'b0;
      end
      if(DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_0_ar_valid) begin
        io_outputs_0_ar_rValid_2 <= 1'b1;
      end
      if(io_outputs_0_ar_validPipe_fire_2) begin
        io_outputs_0_ar_rValid_2 <= 1'b0;
      end
      if(DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_1_ar_valid) begin
        io_outputs_1_ar_rValid_2 <= 1'b1;
      end
      if(io_outputs_1_ar_validPipe_fire_2) begin
        io_outputs_1_ar_rValid_2 <= 1'b0;
      end
      if(DataCachePlugin_setup_dcacheMaster_readOnly_decoder_io_outputs_2_ar_valid) begin
        io_outputs_2_ar_rValid_2 <= 1'b1;
      end
      if(io_outputs_2_ar_validPipe_fire_2) begin
        io_outputs_2_ar_rValid_2 <= 1'b0;
      end
      if(DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_0_aw_valid) begin
        io_outputs_0_aw_rValid_2 <= 1'b1;
      end
      if(io_outputs_0_aw_validPipe_fire_2) begin
        io_outputs_0_aw_rValid_2 <= 1'b0;
      end
      if(DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_1_aw_valid) begin
        io_outputs_1_aw_rValid_2 <= 1'b1;
      end
      if(io_outputs_1_aw_validPipe_fire_2) begin
        io_outputs_1_aw_rValid_2 <= 1'b0;
      end
      if(DataCachePlugin_setup_dcacheMaster_writeOnly_decoder_io_outputs_2_aw_valid) begin
        io_outputs_2_aw_rValid_2 <= 1'b1;
      end
      if(io_outputs_2_aw_validPipe_fire_2) begin
        io_outputs_2_aw_rValid_2 <= 1'b0;
      end
      if(CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_0_ar_valid) begin
        io_outputs_0_ar_rValid_3 <= 1'b1;
      end
      if(io_outputs_0_ar_validPipe_fire_3) begin
        io_outputs_0_ar_rValid_3 <= 1'b0;
      end
      if(CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_1_ar_valid) begin
        io_outputs_1_ar_rValid_3 <= 1'b1;
      end
      if(io_outputs_1_ar_validPipe_fire_3) begin
        io_outputs_1_ar_rValid_3 <= 1'b0;
      end
      if(CoreMemSysPlugin_logic_roMasters_0_readOnly_decoder_io_outputs_2_ar_valid) begin
        io_outputs_2_ar_rValid_3 <= 1'b1;
      end
      if(io_outputs_2_ar_validPipe_fire_3) begin
        io_outputs_2_ar_rValid_3 <= 1'b0;
      end
      if(CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_0_aw_valid) begin
        io_outputs_0_aw_rValid_3 <= 1'b1;
      end
      if(io_outputs_0_aw_validPipe_fire_3) begin
        io_outputs_0_aw_rValid_3 <= 1'b0;
      end
      if(CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_1_aw_valid) begin
        io_outputs_1_aw_rValid_3 <= 1'b1;
      end
      if(io_outputs_1_aw_validPipe_fire_3) begin
        io_outputs_1_aw_rValid_3 <= 1'b0;
      end
      if(CoreMemSysPlugin_logic_roMasters_0_writeOnly_decoder_io_outputs_2_aw_valid) begin
        io_outputs_2_aw_rValid_3 <= 1'b1;
      end
      if(io_outputs_2_aw_validPipe_fire_3) begin
        io_outputs_2_aw_rValid_3 <= 1'b0;
      end
      if(when_CoreNSCSCC_l598) begin
        _zz_io_leds <= (! _zz_io_leds);
      end
    end
  end

  always @(posedge clk) begin
    if(DataCachePlugin_setup_cache_io_mem_read_cmd_ready) begin
      io_mem_read_cmd_rData_id <= DataCachePlugin_setup_cache_io_mem_read_cmd_payload_id;
      io_mem_read_cmd_rData_address <= DataCachePlugin_setup_cache_io_mem_read_cmd_payload_address;
    end
    if(DataCachePlugin_setup_dcacheMaster_r_ready) begin
      DataCachePlugin_setup_dcacheMaster_r_rData_data <= DataCachePlugin_setup_dcacheMaster_r_payload_data;
      DataCachePlugin_setup_dcacheMaster_r_rData_id <= DataCachePlugin_setup_dcacheMaster_r_payload_id;
      DataCachePlugin_setup_dcacheMaster_r_rData_resp <= DataCachePlugin_setup_dcacheMaster_r_payload_resp;
      DataCachePlugin_setup_dcacheMaster_r_rData_last <= DataCachePlugin_setup_dcacheMaster_r_payload_last;
    end
    if(io_mem_toAxi4_awFiltred_ready) begin
      io_mem_toAxi4_awFiltred_rData_last <= io_mem_toAxi4_awFiltred_payload_last;
      io_mem_toAxi4_awFiltred_rData_fragment_address <= io_mem_toAxi4_awFiltred_payload_fragment_address;
      io_mem_toAxi4_awFiltred_rData_fragment_data <= io_mem_toAxi4_awFiltred_payload_fragment_data;
      io_mem_toAxi4_awFiltred_rData_fragment_id <= io_mem_toAxi4_awFiltred_payload_fragment_id;
    end
    if(io_mem_toAxi4_w_ready) begin
      io_mem_toAxi4_w_rData_last <= io_mem_toAxi4_w_payload_last;
      io_mem_toAxi4_w_rData_fragment_address <= io_mem_toAxi4_w_payload_fragment_address;
      io_mem_toAxi4_w_rData_fragment_data <= io_mem_toAxi4_w_payload_fragment_data;
      io_mem_toAxi4_w_rData_fragment_id <= io_mem_toAxi4_w_payload_fragment_id;
    end
    if(DataCachePlugin_setup_dcacheMaster_b_ready) begin
      DataCachePlugin_setup_dcacheMaster_b_rData_id <= DataCachePlugin_setup_dcacheMaster_b_payload_id;
      DataCachePlugin_setup_dcacheMaster_b_rData_resp <= DataCachePlugin_setup_dcacheMaster_b_payload_resp;
    end
    DecodePlugin_logic_debugLA32RDecodedPhysSrc2_idx <= _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_idx;
    DecodePlugin_logic_debugLA32RDecodedPhysSrc2_rtype <= _zz_DecodePlugin_logic_decodedUopsOutputVec_0_archSrc2_rtype;
    DecodePlugin_logic_debugLA32RRawInstruction <= s0_Decode_IssuePipelineSignals_RAW_INSTRUCTIONS_IN_0;
    DispatchPlugin_logic_debugDispatchedUopSrc2_iq0 <= s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
    DispatchPlugin_logic_debugDispatchedUopSrc1_iq0 <= s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
    DispatchPlugin_logic_debugDispatchedUopSrc2_iq1 <= s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
    DispatchPlugin_logic_debugDispatchedUopSrc1_iq1 <= s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
    DispatchPlugin_logic_debugDispatchedUopSrc2_iq2 <= s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
    DispatchPlugin_logic_debugDispatchedUopSrc1_iq2 <= s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
    DispatchPlugin_logic_debugDispatchedUopSrc2_iq3 <= s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
    DispatchPlugin_logic_debugDispatchedUopSrc1_iq3 <= s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
    _zz_io_iqEntryIn_payload_robPtr_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_robPtr;
    _zz_io_iqEntryIn_payload_physDest_idx_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_physDest_idx;
    _zz_io_iqEntryIn_payload_physDestIsFpr_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_physDestIsFpr;
    _zz_io_iqEntryIn_payload_writesToPhysReg_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_writesToPhysReg;
    _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_valid <= AluIntEU_AluIntEuPlugin_euInputPort_payload_useSrc1;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data_2 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Data;
    _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_address <= AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Tag;
    _zz_io_iqEntryIn_payload_src1Ready_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_src1Ready;
    _zz_io_iqEntryIn_payload_src1IsFpr_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_src1IsFpr;
    _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_valid <= AluIntEU_AluIntEuPlugin_euInputPort_payload_useSrc2;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data_2 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Data;
    _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_address <= AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Tag;
    _zz_io_iqEntryIn_payload_src2Ready_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_src2Ready;
    _zz_io_iqEntryIn_payload_src2IsFpr_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_src2IsFpr;
    _zz_io_iqEntryIn_payload_aluCtrl_valid_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_valid;
    _zz_io_iqEntryIn_payload_aluCtrl_isSub_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isSub;
    _zz_io_iqEntryIn_payload_aluCtrl_isAdd_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isAdd;
    _zz_io_iqEntryIn_payload_aluCtrl_isSigned_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_aluCtrl_isSigned;
    _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1 <= _zz_io_iqEntryIn_payload_aluCtrl_logicOp_2;
    _zz_io_iqEntryIn_payload_shiftCtrl_valid_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_valid;
    _zz_io_iqEntryIn_payload_shiftCtrl_isRight_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isRight;
    _zz_io_iqEntryIn_payload_shiftCtrl_isArithmetic_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isArithmetic;
    _zz_io_iqEntryIn_payload_shiftCtrl_isRotate_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isRotate;
    _zz_io_iqEntryIn_payload_shiftCtrl_isDoubleWord_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_shiftCtrl_isDoubleWord;
    _zz_io_iqEntryIn_payload_imm_1 <= AluIntEU_AluIntEuPlugin_euInputPort_payload_imm;
    _zz_io_iqEntryIn_payload_immUsage_1 <= _zz_io_iqEntryIn_payload_immUsage_2;
    _zz_io_iqEntryIn_payload_robPtr <= _zz_io_iqEntryIn_payload_robPtr_1;
    _zz_io_iqEntryIn_payload_physDest_idx <= _zz_io_iqEntryIn_payload_physDest_idx_1;
    _zz_io_iqEntryIn_payload_physDestIsFpr <= _zz_io_iqEntryIn_payload_physDestIsFpr_1;
    _zz_io_iqEntryIn_payload_writesToPhysReg <= _zz_io_iqEntryIn_payload_writesToPhysReg_1;
    _zz_io_iqEntryIn_payload_useSrc1 <= _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_valid;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data_1 <= _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data_2;
    _zz_io_iqEntryIn_payload_src1Tag <= _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_0_address;
    _zz_io_iqEntryIn_payload_src1Ready <= _zz_io_iqEntryIn_payload_src1Ready_1;
    _zz_io_iqEntryIn_payload_src1IsFpr <= _zz_io_iqEntryIn_payload_src1IsFpr_1;
    _zz_io_iqEntryIn_payload_useSrc2 <= _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_valid;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data_1 <= _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data_2;
    _zz_io_iqEntryIn_payload_src2Tag <= _zz_AluIntEU_AluIntEuPlugin_gprReadPorts_1_address;
    _zz_io_iqEntryIn_payload_src2Ready <= _zz_io_iqEntryIn_payload_src2Ready_1;
    _zz_io_iqEntryIn_payload_src2IsFpr <= _zz_io_iqEntryIn_payload_src2IsFpr_1;
    _zz_io_iqEntryIn_payload_aluCtrl_valid <= _zz_io_iqEntryIn_payload_aluCtrl_valid_1;
    _zz_io_iqEntryIn_payload_aluCtrl_isSub <= _zz_io_iqEntryIn_payload_aluCtrl_isSub_1;
    _zz_io_iqEntryIn_payload_aluCtrl_isAdd <= _zz_io_iqEntryIn_payload_aluCtrl_isAdd_1;
    _zz_io_iqEntryIn_payload_aluCtrl_isSigned <= _zz_io_iqEntryIn_payload_aluCtrl_isSigned_1;
    _zz_io_iqEntryIn_payload_aluCtrl_logicOp <= _zz_io_iqEntryIn_payload_aluCtrl_logicOp_1;
    _zz_io_iqEntryIn_payload_shiftCtrl_valid <= _zz_io_iqEntryIn_payload_shiftCtrl_valid_1;
    _zz_io_iqEntryIn_payload_shiftCtrl_isRight <= _zz_io_iqEntryIn_payload_shiftCtrl_isRight_1;
    _zz_io_iqEntryIn_payload_shiftCtrl_isArithmetic <= _zz_io_iqEntryIn_payload_shiftCtrl_isArithmetic_1;
    _zz_io_iqEntryIn_payload_shiftCtrl_isRotate <= _zz_io_iqEntryIn_payload_shiftCtrl_isRotate_1;
    _zz_io_iqEntryIn_payload_shiftCtrl_isDoubleWord <= _zz_io_iqEntryIn_payload_shiftCtrl_isDoubleWord_1;
    _zz_io_iqEntryIn_payload_imm <= _zz_io_iqEntryIn_payload_imm_1;
    _zz_io_iqEntryIn_payload_immUsage <= _zz_io_iqEntryIn_payload_immUsage_1;
    _zz_io_iqEntryIn_payload_src1Data <= AluIntEU_AluIntEuPlugin_gprReadPorts_0_rsp;
    _zz_io_iqEntryIn_payload_src2Data <= AluIntEU_AluIntEuPlugin_gprReadPorts_1_rsp;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_robPtr <= _zz_io_iqEntryIn_payload_robPtr;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_physDest_idx <= _zz_io_iqEntryIn_payload_physDest_idx;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_physDestIsFpr <= _zz_io_iqEntryIn_payload_physDestIsFpr;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_writesToPhysReg <= _zz_io_iqEntryIn_payload_writesToPhysReg;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_useSrc1 <= _zz_io_iqEntryIn_payload_useSrc1;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data <= _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Data_1;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Tag <= _zz_io_iqEntryIn_payload_src1Tag;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1Ready <= _zz_io_iqEntryIn_payload_src1Ready;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src1IsFpr <= _zz_io_iqEntryIn_payload_src1IsFpr;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_useSrc2 <= _zz_io_iqEntryIn_payload_useSrc2;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data <= _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Data_1;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Tag <= _zz_io_iqEntryIn_payload_src2Tag;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2Ready <= _zz_io_iqEntryIn_payload_src2Ready;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_src2IsFpr <= _zz_io_iqEntryIn_payload_src2IsFpr;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_valid <= _zz_io_iqEntryIn_payload_aluCtrl_valid;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSub <= _zz_io_iqEntryIn_payload_aluCtrl_isSub;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isAdd <= _zz_io_iqEntryIn_payload_aluCtrl_isAdd;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_isSigned <= _zz_io_iqEntryIn_payload_aluCtrl_isSigned;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_aluCtrl_logicOp <= _zz_io_iqEntryIn_payload_aluCtrl_logicOp;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_valid <= _zz_io_iqEntryIn_payload_shiftCtrl_valid;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRight <= _zz_io_iqEntryIn_payload_shiftCtrl_isRight;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isArithmetic <= _zz_io_iqEntryIn_payload_shiftCtrl_isArithmetic;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isRotate <= _zz_io_iqEntryIn_payload_shiftCtrl_isRotate;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_shiftCtrl_isDoubleWord <= _zz_io_iqEntryIn_payload_shiftCtrl_isDoubleWord;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_imm <= _zz_io_iqEntryIn_payload_imm;
    _zz_AluIntEU_AluIntEuPlugin_euResult_uop_immUsage <= _zz_io_iqEntryIn_payload_immUsage;
    _zz_AluIntEU_AluIntEuPlugin_euResult_data <= AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_data;
    _zz_AluIntEU_AluIntEuPlugin_euResult_writesToPreg <= AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_writesToPhysReg;
    _zz_AluIntEU_AluIntEuPlugin_euResult_hasException <= AluIntEU_AluIntEuPlugin_intAlu_io_resultOut_payload_hasException;
    _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode <= _zz_AluIntEU_AluIntEuPlugin_euResult_exceptionCode_1;
    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_6 <= MulEU_MulEuPlugin_euInputPort_payload_robPtr;
    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_6 <= MulEU_MulEuPlugin_euInputPort_payload_physDest_idx;
    _zz_MulEU_MulEuPlugin_euResult_writesToPreg_6 <= MulEU_MulEuPlugin_euInputPort_payload_writesToPhysReg;
    _zz_MulEU_MulEuPlugin_gprReadPorts_0_valid <= MulEU_MulEuPlugin_euInputPort_payload_useSrc1;
    _zz_MulEU_MulEuPlugin_gprReadPorts_0_address <= MulEU_MulEuPlugin_euInputPort_payload_src1Tag;
    _zz_MulEU_MulEuPlugin_gprReadPorts_1_valid <= MulEU_MulEuPlugin_euInputPort_payload_useSrc2;
    _zz_MulEU_MulEuPlugin_gprReadPorts_1_address <= MulEU_MulEuPlugin_euInputPort_payload_src2Tag;
    _zz_23 <= MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isDiv;
    _zz_24 <= MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isSigned;
    _zz_25 <= MulEU_MulEuPlugin_euInputPort_payload_mulDivCtrl_isWordOp;
    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_4 <= _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_6;
    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_4 <= _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_6;
    _zz_MulEU_MulEuPlugin_euResult_writesToPreg_4 <= _zz_MulEU_MulEuPlugin_euResult_writesToPreg_6;
    _zz_17 <= _zz_23;
    _zz_18 <= _zz_24;
    _zz_19 <= _zz_25;
    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_3 <= _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_4;
    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_3 <= _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_4;
    _zz_MulEU_MulEuPlugin_euResult_writesToPreg_3 <= _zz_MulEU_MulEuPlugin_euResult_writesToPreg_4;
    _zz_14 <= _zz_17;
    _zz_15 <= _zz_18;
    _zz_16 <= _zz_19;
    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_2 <= _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_3;
    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_2 <= _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_3;
    _zz_MulEU_MulEuPlugin_euResult_writesToPreg_2 <= _zz_MulEU_MulEuPlugin_euResult_writesToPreg_3;
    _zz_11 <= _zz_14;
    _zz_12 <= _zz_15;
    _zz_13 <= _zz_16;
    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_1 <= _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_2;
    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_1 <= _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_2;
    _zz_MulEU_MulEuPlugin_euResult_writesToPreg_1 <= _zz_MulEU_MulEuPlugin_euResult_writesToPreg_2;
    _zz_8 <= _zz_11;
    _zz_9 <= _zz_12;
    _zz_10 <= _zz_13;
    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr <= _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_1;
    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx <= _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_1;
    _zz_MulEU_MulEuPlugin_euResult_writesToPreg <= _zz_MulEU_MulEuPlugin_euResult_writesToPreg_1;
    _zz_5 <= _zz_8;
    _zz_6 <= _zz_9;
    _zz_7 <= _zz_10;
    _zz_MulEU_MulEuPlugin_euResult_uop_robPtr_5 <= _zz_MulEU_MulEuPlugin_euResult_uop_robPtr;
    _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx_5 <= _zz_MulEU_MulEuPlugin_euResult_uop_physDest_idx;
    _zz_MulEU_MulEuPlugin_euResult_writesToPreg_5 <= _zz_MulEU_MulEuPlugin_euResult_writesToPreg;
    _zz_20 <= _zz_5;
    _zz_21 <= _zz_6;
    _zz_22 <= _zz_7;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_robPtr;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_physDest_idx;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_physDestIsFpr;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_writesToPhysReg;
    _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_valid <= BranchEU_BranchEuPlugin_euInputPort_payload_useSrc1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_src1Data;
    _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_address <= BranchEU_BranchEuPlugin_euInputPort_payload_src1Tag;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_src1Ready;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_src1IsFpr;
    _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_valid <= BranchEU_BranchEuPlugin_euInputPort_payload_useSrc2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_src2Data;
    _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_address <= BranchEU_BranchEuPlugin_euInputPort_payload_src2Tag;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_src2Ready;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_src2IsFpr;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_3;
    _zz_switch_BranchEuPlugin_l133 <= BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isJump;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isLink;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_linkReg_idx;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_3;
    _zz_switch_BranchEuPlugin_l133_1 <= BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_isIndirect;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_branchCtrl_laCfIdx;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_imm;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_2 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_3;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_isTaken;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_target;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted_2 <= BranchEU_BranchEuPlugin_euInputPort_payload_branchPrediction_wasPredicted;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc1_1 <= _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_valid;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Tag_1 <= _zz_BranchEU_BranchEuPlugin_gprReadPorts_0_address;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc2_1 <= _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_valid;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Tag_1 <= _zz_BranchEU_BranchEuPlugin_gprReadPorts_1_address;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump_1 <= _zz_switch_BranchEuPlugin_l133;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect_1 <= _zz_switch_BranchEuPlugin_l133_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target_2;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted_1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted_2;
    _zz_BranchEU_BranchEuPlugin_euResult_data_2 <= _zz_BranchEU_BranchEuPlugin_euResult_data_3;
    _zz_BranchEU_BranchEuPlugin_euResult_data_1 <= _zz_BranchEU_BranchEuPlugin_euResult_data_4;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr <= _zz_BranchEU_BranchEuPlugin_euResult_uop_robPtr_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx <= _zz_BranchEU_BranchEuPlugin_euResult_uop_physDest_idx_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr <= _zz_BranchEU_BranchEuPlugin_euResult_uop_physDestIsFpr_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg <= _zz_BranchEU_BranchEuPlugin_euResult_uop_writesToPhysReg_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc1 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc1_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Data_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Tag <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Tag_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src1Ready_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src1IsFpr_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc2 <= _zz_BranchEU_BranchEuPlugin_euResult_uop_useSrc2_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Data_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Tag <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Tag_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src2Ready_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr <= _zz_BranchEU_BranchEuPlugin_euResult_uop_src2IsFpr_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_condition_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isJump_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_idx_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_linkReg_rtype_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isIndirect_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_laCfIdx_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_imm <= _zz_BranchEU_BranchEuPlugin_euResult_uop_imm_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_pc <= _zz_BranchEU_BranchEuPlugin_euResult_uop_pc_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_isTaken_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_target_1;
    _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchPrediction_wasPredicted_1;
    _zz_BranchEU_BranchEuPlugin_euResult_isMispredictedBranch <= (! _zz_BranchEU_BranchEuPlugin_euResult_isMispredictedBranch_1);
    _zz_BranchEU_BranchEuPlugin_euResult_isTaken <= _zz_BranchEU_BranchEuPlugin_euResult_isTaken_1;
    _zz_BranchEU_BranchEuPlugin_euResult_writesToPreg <= _zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink_1;
    _zz_BranchEU_BranchEuPlugin_euResult_data <= (_zz_BranchEU_BranchEuPlugin_euResult_uop_branchCtrl_isLink_1 ? _zz_BranchEU_BranchEuPlugin_euResult_data_5 : _zz_BranchEU_BranchEuPlugin_euResult_data_6);
    if(s0_Decode_ready_output) begin
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_pc <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_pc;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isValid <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isValid;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_uopCode;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_exeUnit;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isa;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1 <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2 <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_imm <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_imm;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_immUsage;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1 <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2 <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1 <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isSerializing <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isSerializing;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target;
      s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted <= s0_Decode_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted;
    end
    if(s1_Rename_ready_output) begin
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_pc <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_pc;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isValid <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isValid;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_uopCode <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_uopCode;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_exeUnit <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_exeUnit;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isa <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isa;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_idx;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archDest_rtype;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_writeArchDestEn;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_idx;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc1_rtype;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1 <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc1;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_idx;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_archSrc2_rtype;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2 <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_useArchSrc2;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_usePcForAddr;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_imm <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_imm;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_immUsage <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_immUsage;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_valid;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSub;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isAdd;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_isSigned;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_aluCtrl_logicOp;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_valid;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRight;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isArithmetic;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isRotate;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_shiftCtrl_isDoubleWord;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_valid;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isDiv;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isSigned;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_mulDivCtrl_isWordOp;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_size;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isSignedLoad;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStore;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isLoadLinked;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isStoreCond;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_atomicOp;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isFence;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_fenceMode;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isCacheOp;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_cacheOpType;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_memCtrl_isPrefetch;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_condition;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isJump;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isLink;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_idx;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_linkReg_rtype;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_isIndirect;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchCtrl_laCfIdx;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_opType;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1 <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc1;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2 <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeSrc2;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fpSizeDest;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_roundingMode;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isIntegerDest;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_isSignedCvt;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1 <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fmaNegSrc1;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_fpuCtrl_fcmpCond;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_csrAddr;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isWrite;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isRead;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_isExchange;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_csrCtrl_useUimmAsSrc;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_sysCode;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isExceptionReturn;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_isTlbOp;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_sysCtrl_tlbOpType;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_decodeExceptionCode;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_hasDecodeException;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isMicrocode;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_microcodeEntry;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isSerializing <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isSerializing;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_isBranchOrJump;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_isTaken;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_target;
      s2_RobAlloc_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted <= s1_Rename_IssuePipelineSignals_DECODED_UOPS_0_branchPrediction_wasPredicted;
      s2_RobAlloc_IssuePipelineSignals_NEEDS_PHYS_REG_0 <= s1_Rename_IssuePipelineSignals_NEEDS_PHYS_REG_0;
    end
    if(s2_RobAlloc_ready_output) begin
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_pc;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isValid;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_uopCode;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_exeUnit;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isa;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_idx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archDest_rtype;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_writeArchDestEn;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_idx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc1_rtype;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1 <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc1;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_idx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_archSrc2_rtype;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2 <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_useArchSrc2;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_usePcForAddr;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_imm;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_immUsage;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_valid;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSub;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isAdd;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_isSigned;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_aluCtrl_logicOp;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_valid;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRight;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isArithmetic;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isRotate;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_shiftCtrl_isDoubleWord;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_valid;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isDiv;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isSigned;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_mulDivCtrl_isWordOp;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_size;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isSignedLoad;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStore;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isLoadLinked;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isStoreCond;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_atomicOp;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isFence;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_fenceMode;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isCacheOp;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_cacheOpType;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_memCtrl_isPrefetch;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_condition;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isJump;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isLink;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_idx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_linkReg_rtype;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_isIndirect;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchCtrl_laCfIdx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_opType;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1 <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc1;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2 <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeSrc2;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fpSizeDest;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_roundingMode;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isIntegerDest;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_isSignedCvt;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1 <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fmaNegSrc1;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_fpuCtrl_fcmpCond;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_csrAddr;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isWrite;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isRead;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_isExchange;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_csrCtrl_useUimmAsSrc;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_sysCode;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isExceptionReturn;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_isTlbOp;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_sysCtrl_tlbOpType;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_decodeExceptionCode;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_hasDecodeException;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isMicrocode;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_microcodeEntry;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isSerializing;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_isBranchOrJump;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_isTaken;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_target;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_decoded_branchPrediction_wasPredicted;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1_idx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc1IsFpr;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2_idx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physSrc2IsFpr;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDest_idx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_physDestIsFpr;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDest_idx;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_oldPhysDestIsFpr;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_allocatesPhysDest;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_rename_writesToPhysReg;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_robPtr;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_uniqueId;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_dispatched;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_executed <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_executed;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_hasException;
      s3_Dispatch_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode <= s2_RobAlloc_IssuePipelineSignals_ALLOCATED_UOPS_0_exceptionCode;
    end
    if(_zz_LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_valid) begin
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_qPtr;
      _zz_when_AddressGenerationUnit_l215 <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_basePhysReg;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_immediate;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_accessSize;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_usePc;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_pc;
      _zz_when_AddressGenerationUnit_l220 <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_dataReg;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_robPtr;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isLoad;
      _zz_when_AddressGenerationUnit_l220_1 <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isStore;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isFlush;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_isIO;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst <= LsuEU_LsuEuPlugin_hw_aguPort_input_payload_physDst;
    end
    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address <= LsuEU_LsuEuPlugin_hw_aguPort_prfReadBase_rsp;
    _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData <= LsuEU_LsuEuPlugin_hw_aguPort_prfReadData_rsp;
    if(_zz_LsuEU_LsuEuPlugin_hw_aguPort_input_ready) begin
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr_1 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_qPtr;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_5 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_4;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_2 <= (((_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_4 & _zz__zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException_2) != 32'h0) && (_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_alignException != MemAccessSize_B));
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize_2 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_accessSize;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_2 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeMask_1;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_basePhysReg <= _zz_when_AddressGenerationUnit_l215;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate_1 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_immediate;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc_1 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_usePc;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc_1 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_pc;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr_1 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_robPtr;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad_1 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isLoad;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isStore <= _zz_when_AddressGenerationUnit_l220_1;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst_1 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_physDst;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_4 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_storeData_3;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush_1 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isFlush;
      _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO_1 <= (_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_isIO || (1'b0 || ((32'hbfd00000 <= _zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_4) && (_zz_LsuEU_LsuEuPlugin_hw_aguPort_output_payload_address_4 <= 32'hc0100000))));
    end
    if(StoreBufferPlugin_hw_sqQueryPort_cmd_valid) begin
      LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_hit <= StoreBufferPlugin_hw_sqQueryPort_rsp_hit;
      LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_data <= StoreBufferPlugin_hw_sqQueryPort_rsp_data;
      LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_olderStoreHasUnknownAddress <= StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreHasUnknownAddress;
      LoadQueuePlugin_logic_loadQueue_sbQueryRspReg_olderStoreDataNotReady <= StoreBufferPlugin_hw_sqQueryPort_rsp_olderStoreDataNotReady;
    end
    LoadQueuePlugin_logic_loadQueue_completingHead_valid <= LoadQueuePlugin_logic_loadQueue_slots_0_valid;
    LoadQueuePlugin_logic_loadQueue_completingHead_address <= LoadQueuePlugin_logic_loadQueue_slots_0_address;
    LoadQueuePlugin_logic_loadQueue_completingHead_size <= LoadQueuePlugin_logic_loadQueue_slots_0_size;
    LoadQueuePlugin_logic_loadQueue_completingHead_robPtr <= LoadQueuePlugin_logic_loadQueue_slots_0_robPtr;
    LoadQueuePlugin_logic_loadQueue_completingHead_pdest <= LoadQueuePlugin_logic_loadQueue_slots_0_pdest;
    LoadQueuePlugin_logic_loadQueue_completingHead_isIO <= LoadQueuePlugin_logic_loadQueue_slots_0_isIO;
    LoadQueuePlugin_logic_loadQueue_completingHead_hasException <= LoadQueuePlugin_logic_loadQueue_slots_0_hasException;
    LoadQueuePlugin_logic_loadQueue_completingHead_exceptionCode <= LoadQueuePlugin_logic_loadQueue_slots_0_exceptionCode;
    LoadQueuePlugin_logic_loadQueue_completingHead_isWaitingForFwdRsp <= LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForFwdRsp;
    LoadQueuePlugin_logic_loadQueue_completingHead_isStalledByDependency <= LoadQueuePlugin_logic_loadQueue_slots_0_isStalledByDependency;
    LoadQueuePlugin_logic_loadQueue_completingHead_isReadyForDCache <= LoadQueuePlugin_logic_loadQueue_slots_0_isReadyForDCache;
    LoadQueuePlugin_logic_loadQueue_completingHead_isWaitingForRsp <= LoadQueuePlugin_logic_loadQueue_slots_0_isWaitingForRsp;
    if(s1_PC_Gen_ready_output) begin
      s2_ICache_Access_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC <= s1_PC_Gen_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC;
      s2_ICache_Access_FetchPipelinePlugin_logic_FetchPipeline_PC <= s1_PC_Gen_FetchPipelinePlugin_logic_FetchPipeline_PC;
    end
    if(s2_ICache_Access_ready_output) begin
      s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_PC <= s2_ICache_Access_FetchPipelinePlugin_logic_FetchPipeline_PC;
      s4_Predecode_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC <= s2_ICache_Access_FetchPipelinePlugin_logic_FetchPipeline_RAW_PC;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_IDLE_OH_ID]) : begin
        if(when_ICachePlugin_l212) begin
          ICachePlugin_logic_refill_refillCmdReg_address <= ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_address;
          ICachePlugin_logic_refill_refillCmdReg_transactionId <= ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_transactionId;
          ICachePlugin_logic_refill_victimWayReg <= ICachePlugin_logic_pipeline_f2_f2_metaLine_lru;
          ICachePlugin_logic_refill_latchedMetaOnMiss_ways_0_tag <= ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_0_tag;
          ICachePlugin_logic_refill_latchedMetaOnMiss_ways_1_tag <= ICachePlugin_logic_pipeline_f2_f2_metaLine_ways_1_tag;
          ICachePlugin_logic_refill_latchedMetaOnMiss_lru <= ICachePlugin_logic_pipeline_f2_f2_metaLine_lru;
        end
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_SEND_REQ_OH_ID]) : begin
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_RECEIVE_DATA_OH_ID]) : begin
        if(ICachePlugin_axiMaster_r_fire) begin
          if(_zz_78[0]) begin
            ICachePlugin_logic_refill_lineBuffer_0 <= ICachePlugin_axiMaster_r_payload_data;
          end
          if(_zz_78[1]) begin
            ICachePlugin_logic_refill_lineBuffer_1 <= ICachePlugin_axiMaster_r_payload_data;
          end
          if(_zz_78[2]) begin
            ICachePlugin_logic_refill_lineBuffer_2 <= ICachePlugin_axiMaster_r_payload_data;
          end
          if(_zz_78[3]) begin
            ICachePlugin_logic_refill_lineBuffer_3 <= ICachePlugin_axiMaster_r_payload_data;
          end
        end
      end
      (ICachePlugin_logic_refill_fsm_stateReg[ICachePlugin_logic_refill_fsm_COMMIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_address <= ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_address;
    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_CMD_transactionId <= ICache_F1_Access_ICachePlugin_logic_pipeline_F1_CMD_transactionId;
    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_VALID_MASK_0 <= ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_0;
    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F1_VALID_MASK_1 <= ICache_F1_Access_ICachePlugin_logic_pipeline_F1_VALID_MASK_1;
    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_USE_FORWARDED_META <= ICache_F1_Access_ICachePlugin_logic_pipeline_F2_USE_FORWARDED_META;
    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_0_tag <= ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_0_tag;
    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_1_tag <= ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_ways_1_tag;
    ICache_F2_HitCheck_ICachePlugin_logic_pipeline_F2_FORWARDED_META_lru <= ICache_F1_Access_ICachePlugin_logic_pipeline_F2_FORWARDED_META_lru;
    BpuPipelinePlugin_logic_s2_predict_Q_PC <= BpuPipelinePlugin_logic_s1_read_Q_PC;
    BpuPipelinePlugin_logic_s2_predict_TRANSACTION_ID <= BpuPipelinePlugin_logic_s1_read_TRANSACTION_ID;
    BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_pc <= BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_pc;
    BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_isTaken <= BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_isTaken;
    BpuPipelinePlugin_logic_u2_write_U_PAYLOAD_target <= BpuPipelinePlugin_logic_u1_read_U_PAYLOAD_target;
    _zz_when_CoreNSCSCC_l598_1 <= _zz_when_CoreNSCSCC_l598;
  end

  always @(posedge clk) begin
    BpuPipelinePlugin_queryPortIn_payload_pc_regNext <= BpuPipelinePlugin_queryPortIn_payload_pc;
    BpuPipelinePlugin_queryPortIn_payload_transactionId_regNext <= BpuPipelinePlugin_queryPortIn_payload_transactionId;
  end


endmodule

module BufferCC (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          clk,
  input  wire          reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk) begin
    buffers_0 <= io_dataIn;
    buffers_1 <= buffers_0;
  end


endmodule

//Axi4WriteOnlyArbiter_2 replaced by Axi4WriteOnlyArbiter

//Axi4ReadOnlyArbiter_2 replaced by Axi4ReadOnlyArbiter

//Axi4WriteOnlyArbiter_1 replaced by Axi4WriteOnlyArbiter

//Axi4ReadOnlyArbiter_1 replaced by Axi4ReadOnlyArbiter

module Axi4WriteOnlyArbiter (
  input  wire          io_inputs_0_aw_valid,
  output wire          io_inputs_0_aw_ready,
  input  wire [31:0]   io_inputs_0_aw_payload_addr,
  input  wire [4:0]    io_inputs_0_aw_payload_id,
  input  wire [7:0]    io_inputs_0_aw_payload_len,
  input  wire [2:0]    io_inputs_0_aw_payload_size,
  input  wire [1:0]    io_inputs_0_aw_payload_burst,
  input  wire          io_inputs_0_w_valid,
  output wire          io_inputs_0_w_ready,
  input  wire [31:0]   io_inputs_0_w_payload_data,
  input  wire [3:0]    io_inputs_0_w_payload_strb,
  input  wire          io_inputs_0_w_payload_last,
  output wire          io_inputs_0_b_valid,
  input  wire          io_inputs_0_b_ready,
  output wire [4:0]    io_inputs_0_b_payload_id,
  output wire [1:0]    io_inputs_0_b_payload_resp,
  input  wire          io_inputs_1_aw_valid,
  output wire          io_inputs_1_aw_ready,
  input  wire [31:0]   io_inputs_1_aw_payload_addr,
  input  wire [4:0]    io_inputs_1_aw_payload_id,
  input  wire [7:0]    io_inputs_1_aw_payload_len,
  input  wire [2:0]    io_inputs_1_aw_payload_size,
  input  wire [1:0]    io_inputs_1_aw_payload_burst,
  input  wire          io_inputs_1_w_valid,
  output wire          io_inputs_1_w_ready,
  input  wire [31:0]   io_inputs_1_w_payload_data,
  input  wire [3:0]    io_inputs_1_w_payload_strb,
  input  wire          io_inputs_1_w_payload_last,
  output wire          io_inputs_1_b_valid,
  input  wire          io_inputs_1_b_ready,
  output wire [4:0]    io_inputs_1_b_payload_id,
  output wire [1:0]    io_inputs_1_b_payload_resp,
  input  wire          io_inputs_2_aw_valid,
  output wire          io_inputs_2_aw_ready,
  input  wire [31:0]   io_inputs_2_aw_payload_addr,
  input  wire [4:0]    io_inputs_2_aw_payload_id,
  input  wire [7:0]    io_inputs_2_aw_payload_len,
  input  wire [2:0]    io_inputs_2_aw_payload_size,
  input  wire [1:0]    io_inputs_2_aw_payload_burst,
  input  wire          io_inputs_2_w_valid,
  output wire          io_inputs_2_w_ready,
  input  wire [31:0]   io_inputs_2_w_payload_data,
  input  wire [3:0]    io_inputs_2_w_payload_strb,
  input  wire          io_inputs_2_w_payload_last,
  output wire          io_inputs_2_b_valid,
  input  wire          io_inputs_2_b_ready,
  output wire [4:0]    io_inputs_2_b_payload_id,
  output wire [1:0]    io_inputs_2_b_payload_resp,
  input  wire          io_inputs_3_aw_valid,
  output wire          io_inputs_3_aw_ready,
  input  wire [31:0]   io_inputs_3_aw_payload_addr,
  input  wire [4:0]    io_inputs_3_aw_payload_id,
  input  wire [7:0]    io_inputs_3_aw_payload_len,
  input  wire [2:0]    io_inputs_3_aw_payload_size,
  input  wire [1:0]    io_inputs_3_aw_payload_burst,
  input  wire          io_inputs_3_w_valid,
  output wire          io_inputs_3_w_ready,
  input  wire [31:0]   io_inputs_3_w_payload_data,
  input  wire [3:0]    io_inputs_3_w_payload_strb,
  input  wire          io_inputs_3_w_payload_last,
  output wire          io_inputs_3_b_valid,
  input  wire          io_inputs_3_b_ready,
  output wire [4:0]    io_inputs_3_b_payload_id,
  output wire [1:0]    io_inputs_3_b_payload_resp,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [6:0]    io_output_aw_payload_id,
  output wire [7:0]    io_output_aw_payload_len,
  output wire [2:0]    io_output_aw_payload_size,
  output wire [1:0]    io_output_aw_payload_burst,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [31:0]   io_output_w_payload_data,
  output wire [3:0]    io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [6:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          clk,
  input  wire          reset
);

  reg                 cmdArbiter_io_output_ready;
  wire                cmdRouteFork_translated_fifo_io_pop_ready;
  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_inputs_2_ready;
  wire                cmdArbiter_io_inputs_3_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [31:0]   cmdArbiter_io_output_payload_addr;
  wire       [4:0]    cmdArbiter_io_output_payload_id;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire       [1:0]    cmdArbiter_io_chosen;
  wire       [3:0]    cmdArbiter_io_chosenOH;
  wire                cmdRouteFork_translated_fifo_io_push_ready;
  wire                cmdRouteFork_translated_fifo_io_pop_valid;
  wire       [1:0]    cmdRouteFork_translated_fifo_io_pop_payload;
  wire       [2:0]    cmdRouteFork_translated_fifo_io_occupancy;
  wire       [2:0]    cmdRouteFork_translated_fifo_io_availability;
  reg                 _zz_io_output_w_valid;
  reg        [31:0]   _zz_io_output_w_payload_data;
  reg        [3:0]    _zz_io_output_w_payload_strb;
  reg                 _zz_io_output_w_payload_last;
  reg                 _zz_io_output_b_ready;
  wire                cmdOutputFork_valid;
  wire                cmdOutputFork_ready;
  wire       [31:0]   cmdOutputFork_payload_addr;
  wire       [4:0]    cmdOutputFork_payload_id;
  wire       [7:0]    cmdOutputFork_payload_len;
  wire       [2:0]    cmdOutputFork_payload_size;
  wire       [1:0]    cmdOutputFork_payload_burst;
  wire                cmdRouteFork_valid;
  wire                cmdRouteFork_ready;
  wire       [31:0]   cmdRouteFork_payload_addr;
  wire       [4:0]    cmdRouteFork_payload_id;
  wire       [7:0]    cmdRouteFork_payload_len;
  wire       [2:0]    cmdRouteFork_payload_size;
  wire       [1:0]    cmdRouteFork_payload_burst;
  reg                 cmdArbiter_io_output_fork2_logic_linkEnable_0;
  reg                 cmdArbiter_io_output_fork2_logic_linkEnable_1;
  wire                when_Stream_l1253;
  wire                when_Stream_l1253_1;
  wire                cmdOutputFork_fire;
  wire                cmdRouteFork_fire;
  wire                cmdRouteFork_translated_valid;
  wire                cmdRouteFork_translated_ready;
  wire       [1:0]    cmdRouteFork_translated_payload;
  wire                io_output_w_fire;
  wire       [1:0]    writeRspIndex;
  wire                writeRspSels_0;
  wire                writeRspSels_1;
  wire                writeRspSels_2;
  wire                writeRspSels_3;

  StreamArbiter cmdArbiter (
    .io_inputs_0_valid         (io_inputs_0_aw_valid                   ), //i
    .io_inputs_0_ready         (cmdArbiter_io_inputs_0_ready           ), //o
    .io_inputs_0_payload_addr  (io_inputs_0_aw_payload_addr[31:0]      ), //i
    .io_inputs_0_payload_id    (io_inputs_0_aw_payload_id[4:0]         ), //i
    .io_inputs_0_payload_len   (io_inputs_0_aw_payload_len[7:0]        ), //i
    .io_inputs_0_payload_size  (io_inputs_0_aw_payload_size[2:0]       ), //i
    .io_inputs_0_payload_burst (io_inputs_0_aw_payload_burst[1:0]      ), //i
    .io_inputs_1_valid         (io_inputs_1_aw_valid                   ), //i
    .io_inputs_1_ready         (cmdArbiter_io_inputs_1_ready           ), //o
    .io_inputs_1_payload_addr  (io_inputs_1_aw_payload_addr[31:0]      ), //i
    .io_inputs_1_payload_id    (io_inputs_1_aw_payload_id[4:0]         ), //i
    .io_inputs_1_payload_len   (io_inputs_1_aw_payload_len[7:0]        ), //i
    .io_inputs_1_payload_size  (io_inputs_1_aw_payload_size[2:0]       ), //i
    .io_inputs_1_payload_burst (io_inputs_1_aw_payload_burst[1:0]      ), //i
    .io_inputs_2_valid         (io_inputs_2_aw_valid                   ), //i
    .io_inputs_2_ready         (cmdArbiter_io_inputs_2_ready           ), //o
    .io_inputs_2_payload_addr  (io_inputs_2_aw_payload_addr[31:0]      ), //i
    .io_inputs_2_payload_id    (io_inputs_2_aw_payload_id[4:0]         ), //i
    .io_inputs_2_payload_len   (io_inputs_2_aw_payload_len[7:0]        ), //i
    .io_inputs_2_payload_size  (io_inputs_2_aw_payload_size[2:0]       ), //i
    .io_inputs_2_payload_burst (io_inputs_2_aw_payload_burst[1:0]      ), //i
    .io_inputs_3_valid         (io_inputs_3_aw_valid                   ), //i
    .io_inputs_3_ready         (cmdArbiter_io_inputs_3_ready           ), //o
    .io_inputs_3_payload_addr  (io_inputs_3_aw_payload_addr[31:0]      ), //i
    .io_inputs_3_payload_id    (io_inputs_3_aw_payload_id[4:0]         ), //i
    .io_inputs_3_payload_len   (io_inputs_3_aw_payload_len[7:0]        ), //i
    .io_inputs_3_payload_size  (io_inputs_3_aw_payload_size[2:0]       ), //i
    .io_inputs_3_payload_burst (io_inputs_3_aw_payload_burst[1:0]      ), //i
    .io_output_valid           (cmdArbiter_io_output_valid             ), //o
    .io_output_ready           (cmdArbiter_io_output_ready             ), //i
    .io_output_payload_addr    (cmdArbiter_io_output_payload_addr[31:0]), //o
    .io_output_payload_id      (cmdArbiter_io_output_payload_id[4:0]   ), //o
    .io_output_payload_len     (cmdArbiter_io_output_payload_len[7:0]  ), //o
    .io_output_payload_size    (cmdArbiter_io_output_payload_size[2:0] ), //o
    .io_output_payload_burst   (cmdArbiter_io_output_payload_burst[1:0]), //o
    .io_chosen                 (cmdArbiter_io_chosen[1:0]              ), //o
    .io_chosenOH               (cmdArbiter_io_chosenOH[3:0]            ), //o
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  StreamFifoLowLatency cmdRouteFork_translated_fifo (
    .io_push_valid   (cmdRouteFork_translated_valid                    ), //i
    .io_push_ready   (cmdRouteFork_translated_fifo_io_push_ready       ), //o
    .io_push_payload (cmdRouteFork_translated_payload[1:0]             ), //i
    .io_pop_valid    (cmdRouteFork_translated_fifo_io_pop_valid        ), //o
    .io_pop_ready    (cmdRouteFork_translated_fifo_io_pop_ready        ), //i
    .io_pop_payload  (cmdRouteFork_translated_fifo_io_pop_payload[1:0] ), //o
    .io_flush        (1'b0                                             ), //i
    .io_occupancy    (cmdRouteFork_translated_fifo_io_occupancy[2:0]   ), //o
    .io_availability (cmdRouteFork_translated_fifo_io_availability[2:0]), //o
    .clk             (clk                                              ), //i
    .reset           (reset                                            )  //i
  );
  always @(*) begin
    case(cmdRouteFork_translated_fifo_io_pop_payload)
      2'b00 : begin
        _zz_io_output_w_valid = io_inputs_0_w_valid;
        _zz_io_output_w_payload_data = io_inputs_0_w_payload_data;
        _zz_io_output_w_payload_strb = io_inputs_0_w_payload_strb;
        _zz_io_output_w_payload_last = io_inputs_0_w_payload_last;
      end
      2'b01 : begin
        _zz_io_output_w_valid = io_inputs_1_w_valid;
        _zz_io_output_w_payload_data = io_inputs_1_w_payload_data;
        _zz_io_output_w_payload_strb = io_inputs_1_w_payload_strb;
        _zz_io_output_w_payload_last = io_inputs_1_w_payload_last;
      end
      2'b10 : begin
        _zz_io_output_w_valid = io_inputs_2_w_valid;
        _zz_io_output_w_payload_data = io_inputs_2_w_payload_data;
        _zz_io_output_w_payload_strb = io_inputs_2_w_payload_strb;
        _zz_io_output_w_payload_last = io_inputs_2_w_payload_last;
      end
      default : begin
        _zz_io_output_w_valid = io_inputs_3_w_valid;
        _zz_io_output_w_payload_data = io_inputs_3_w_payload_data;
        _zz_io_output_w_payload_strb = io_inputs_3_w_payload_strb;
        _zz_io_output_w_payload_last = io_inputs_3_w_payload_last;
      end
    endcase
  end

  always @(*) begin
    case(writeRspIndex)
      2'b00 : _zz_io_output_b_ready = io_inputs_0_b_ready;
      2'b01 : _zz_io_output_b_ready = io_inputs_1_b_ready;
      2'b10 : _zz_io_output_b_ready = io_inputs_2_b_ready;
      default : _zz_io_output_b_ready = io_inputs_3_b_ready;
    endcase
  end

  assign io_inputs_0_aw_ready = cmdArbiter_io_inputs_0_ready;
  assign io_inputs_1_aw_ready = cmdArbiter_io_inputs_1_ready;
  assign io_inputs_2_aw_ready = cmdArbiter_io_inputs_2_ready;
  assign io_inputs_3_aw_ready = cmdArbiter_io_inputs_3_ready;
  always @(*) begin
    cmdArbiter_io_output_ready = 1'b1;
    if(when_Stream_l1253) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
    if(when_Stream_l1253_1) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
  end

  assign when_Stream_l1253 = ((! cmdOutputFork_ready) && cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign when_Stream_l1253_1 = ((! cmdRouteFork_ready) && cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdOutputFork_valid = (cmdArbiter_io_output_valid && cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign cmdOutputFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdOutputFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdOutputFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdOutputFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdOutputFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdOutputFork_fire = (cmdOutputFork_valid && cmdOutputFork_ready);
  assign cmdRouteFork_valid = (cmdArbiter_io_output_valid && cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdRouteFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdRouteFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdRouteFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdRouteFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdRouteFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdRouteFork_fire = (cmdRouteFork_valid && cmdRouteFork_ready);
  assign io_output_aw_valid = cmdOutputFork_valid;
  assign cmdOutputFork_ready = io_output_aw_ready;
  assign io_output_aw_payload_addr = cmdOutputFork_payload_addr;
  assign io_output_aw_payload_len = cmdOutputFork_payload_len;
  assign io_output_aw_payload_size = cmdOutputFork_payload_size;
  assign io_output_aw_payload_burst = cmdOutputFork_payload_burst;
  assign io_output_aw_payload_id = {cmdArbiter_io_chosen,cmdArbiter_io_output_payload_id};
  assign cmdRouteFork_translated_valid = cmdRouteFork_valid;
  assign cmdRouteFork_ready = cmdRouteFork_translated_ready;
  assign cmdRouteFork_translated_payload = cmdArbiter_io_chosen;
  assign cmdRouteFork_translated_ready = cmdRouteFork_translated_fifo_io_push_ready;
  assign io_output_w_valid = (cmdRouteFork_translated_fifo_io_pop_valid && _zz_io_output_w_valid);
  assign io_output_w_payload_data = _zz_io_output_w_payload_data;
  assign io_output_w_payload_strb = _zz_io_output_w_payload_strb;
  assign io_output_w_payload_last = _zz_io_output_w_payload_last;
  assign io_inputs_0_w_ready = ((cmdRouteFork_translated_fifo_io_pop_valid && io_output_w_ready) && (cmdRouteFork_translated_fifo_io_pop_payload == 2'b00));
  assign io_inputs_1_w_ready = ((cmdRouteFork_translated_fifo_io_pop_valid && io_output_w_ready) && (cmdRouteFork_translated_fifo_io_pop_payload == 2'b01));
  assign io_inputs_2_w_ready = ((cmdRouteFork_translated_fifo_io_pop_valid && io_output_w_ready) && (cmdRouteFork_translated_fifo_io_pop_payload == 2'b10));
  assign io_inputs_3_w_ready = ((cmdRouteFork_translated_fifo_io_pop_valid && io_output_w_ready) && (cmdRouteFork_translated_fifo_io_pop_payload == 2'b11));
  assign io_output_w_fire = (io_output_w_valid && io_output_w_ready);
  assign cmdRouteFork_translated_fifo_io_pop_ready = (io_output_w_fire && io_output_w_payload_last);
  assign writeRspIndex = io_output_b_payload_id[6 : 5];
  assign writeRspSels_0 = (writeRspIndex == 2'b00);
  assign writeRspSels_1 = (writeRspIndex == 2'b01);
  assign writeRspSels_2 = (writeRspIndex == 2'b10);
  assign writeRspSels_3 = (writeRspIndex == 2'b11);
  assign io_inputs_0_b_valid = (io_output_b_valid && writeRspSels_0);
  assign io_inputs_0_b_payload_resp = io_output_b_payload_resp;
  assign io_inputs_0_b_payload_id = io_output_b_payload_id[4 : 0];
  assign io_inputs_1_b_valid = (io_output_b_valid && writeRspSels_1);
  assign io_inputs_1_b_payload_resp = io_output_b_payload_resp;
  assign io_inputs_1_b_payload_id = io_output_b_payload_id[4 : 0];
  assign io_inputs_2_b_valid = (io_output_b_valid && writeRspSels_2);
  assign io_inputs_2_b_payload_resp = io_output_b_payload_resp;
  assign io_inputs_2_b_payload_id = io_output_b_payload_id[4 : 0];
  assign io_inputs_3_b_valid = (io_output_b_valid && writeRspSels_3);
  assign io_inputs_3_b_payload_resp = io_output_b_payload_resp;
  assign io_inputs_3_b_payload_id = io_output_b_payload_id[4 : 0];
  assign io_output_b_ready = _zz_io_output_b_ready;
  always @(posedge clk) begin
    if(reset) begin
      cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
      cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
    end else begin
      if(cmdOutputFork_fire) begin
        cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdRouteFork_fire) begin
        cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(cmdArbiter_io_output_ready) begin
        cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
        cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
      end
    end
  end


endmodule

module Axi4ReadOnlyArbiter (
  input  wire          io_inputs_0_ar_valid,
  output wire          io_inputs_0_ar_ready,
  input  wire [31:0]   io_inputs_0_ar_payload_addr,
  input  wire [4:0]    io_inputs_0_ar_payload_id,
  input  wire [7:0]    io_inputs_0_ar_payload_len,
  input  wire [2:0]    io_inputs_0_ar_payload_size,
  input  wire [1:0]    io_inputs_0_ar_payload_burst,
  output wire          io_inputs_0_r_valid,
  input  wire          io_inputs_0_r_ready,
  output wire [31:0]   io_inputs_0_r_payload_data,
  output wire [4:0]    io_inputs_0_r_payload_id,
  output wire [1:0]    io_inputs_0_r_payload_resp,
  output wire          io_inputs_0_r_payload_last,
  input  wire          io_inputs_1_ar_valid,
  output wire          io_inputs_1_ar_ready,
  input  wire [31:0]   io_inputs_1_ar_payload_addr,
  input  wire [4:0]    io_inputs_1_ar_payload_id,
  input  wire [7:0]    io_inputs_1_ar_payload_len,
  input  wire [2:0]    io_inputs_1_ar_payload_size,
  input  wire [1:0]    io_inputs_1_ar_payload_burst,
  output wire          io_inputs_1_r_valid,
  input  wire          io_inputs_1_r_ready,
  output wire [31:0]   io_inputs_1_r_payload_data,
  output wire [4:0]    io_inputs_1_r_payload_id,
  output wire [1:0]    io_inputs_1_r_payload_resp,
  output wire          io_inputs_1_r_payload_last,
  input  wire          io_inputs_2_ar_valid,
  output wire          io_inputs_2_ar_ready,
  input  wire [31:0]   io_inputs_2_ar_payload_addr,
  input  wire [4:0]    io_inputs_2_ar_payload_id,
  input  wire [7:0]    io_inputs_2_ar_payload_len,
  input  wire [2:0]    io_inputs_2_ar_payload_size,
  input  wire [1:0]    io_inputs_2_ar_payload_burst,
  output wire          io_inputs_2_r_valid,
  input  wire          io_inputs_2_r_ready,
  output wire [31:0]   io_inputs_2_r_payload_data,
  output wire [4:0]    io_inputs_2_r_payload_id,
  output wire [1:0]    io_inputs_2_r_payload_resp,
  output wire          io_inputs_2_r_payload_last,
  input  wire          io_inputs_3_ar_valid,
  output wire          io_inputs_3_ar_ready,
  input  wire [31:0]   io_inputs_3_ar_payload_addr,
  input  wire [4:0]    io_inputs_3_ar_payload_id,
  input  wire [7:0]    io_inputs_3_ar_payload_len,
  input  wire [2:0]    io_inputs_3_ar_payload_size,
  input  wire [1:0]    io_inputs_3_ar_payload_burst,
  output wire          io_inputs_3_r_valid,
  input  wire          io_inputs_3_r_ready,
  output wire [31:0]   io_inputs_3_r_payload_data,
  output wire [4:0]    io_inputs_3_r_payload_id,
  output wire [1:0]    io_inputs_3_r_payload_resp,
  output wire          io_inputs_3_r_payload_last,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [6:0]    io_output_ar_payload_id,
  output wire [7:0]    io_output_ar_payload_len,
  output wire [2:0]    io_output_ar_payload_size,
  output wire [1:0]    io_output_ar_payload_burst,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [31:0]   io_output_r_payload_data,
  input  wire [6:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_inputs_2_ready;
  wire                cmdArbiter_io_inputs_3_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [31:0]   cmdArbiter_io_output_payload_addr;
  wire       [4:0]    cmdArbiter_io_output_payload_id;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire       [1:0]    cmdArbiter_io_chosen;
  wire       [3:0]    cmdArbiter_io_chosenOH;
  reg                 _zz_io_output_r_ready;
  wire       [1:0]    readRspIndex;
  wire                readRspSels_0;
  wire                readRspSels_1;
  wire                readRspSels_2;
  wire                readRspSels_3;

  StreamArbiter cmdArbiter (
    .io_inputs_0_valid         (io_inputs_0_ar_valid                   ), //i
    .io_inputs_0_ready         (cmdArbiter_io_inputs_0_ready           ), //o
    .io_inputs_0_payload_addr  (io_inputs_0_ar_payload_addr[31:0]      ), //i
    .io_inputs_0_payload_id    (io_inputs_0_ar_payload_id[4:0]         ), //i
    .io_inputs_0_payload_len   (io_inputs_0_ar_payload_len[7:0]        ), //i
    .io_inputs_0_payload_size  (io_inputs_0_ar_payload_size[2:0]       ), //i
    .io_inputs_0_payload_burst (io_inputs_0_ar_payload_burst[1:0]      ), //i
    .io_inputs_1_valid         (io_inputs_1_ar_valid                   ), //i
    .io_inputs_1_ready         (cmdArbiter_io_inputs_1_ready           ), //o
    .io_inputs_1_payload_addr  (io_inputs_1_ar_payload_addr[31:0]      ), //i
    .io_inputs_1_payload_id    (io_inputs_1_ar_payload_id[4:0]         ), //i
    .io_inputs_1_payload_len   (io_inputs_1_ar_payload_len[7:0]        ), //i
    .io_inputs_1_payload_size  (io_inputs_1_ar_payload_size[2:0]       ), //i
    .io_inputs_1_payload_burst (io_inputs_1_ar_payload_burst[1:0]      ), //i
    .io_inputs_2_valid         (io_inputs_2_ar_valid                   ), //i
    .io_inputs_2_ready         (cmdArbiter_io_inputs_2_ready           ), //o
    .io_inputs_2_payload_addr  (io_inputs_2_ar_payload_addr[31:0]      ), //i
    .io_inputs_2_payload_id    (io_inputs_2_ar_payload_id[4:0]         ), //i
    .io_inputs_2_payload_len   (io_inputs_2_ar_payload_len[7:0]        ), //i
    .io_inputs_2_payload_size  (io_inputs_2_ar_payload_size[2:0]       ), //i
    .io_inputs_2_payload_burst (io_inputs_2_ar_payload_burst[1:0]      ), //i
    .io_inputs_3_valid         (io_inputs_3_ar_valid                   ), //i
    .io_inputs_3_ready         (cmdArbiter_io_inputs_3_ready           ), //o
    .io_inputs_3_payload_addr  (io_inputs_3_ar_payload_addr[31:0]      ), //i
    .io_inputs_3_payload_id    (io_inputs_3_ar_payload_id[4:0]         ), //i
    .io_inputs_3_payload_len   (io_inputs_3_ar_payload_len[7:0]        ), //i
    .io_inputs_3_payload_size  (io_inputs_3_ar_payload_size[2:0]       ), //i
    .io_inputs_3_payload_burst (io_inputs_3_ar_payload_burst[1:0]      ), //i
    .io_output_valid           (cmdArbiter_io_output_valid             ), //o
    .io_output_ready           (io_output_ar_ready                     ), //i
    .io_output_payload_addr    (cmdArbiter_io_output_payload_addr[31:0]), //o
    .io_output_payload_id      (cmdArbiter_io_output_payload_id[4:0]   ), //o
    .io_output_payload_len     (cmdArbiter_io_output_payload_len[7:0]  ), //o
    .io_output_payload_size    (cmdArbiter_io_output_payload_size[2:0] ), //o
    .io_output_payload_burst   (cmdArbiter_io_output_payload_burst[1:0]), //o
    .io_chosen                 (cmdArbiter_io_chosen[1:0]              ), //o
    .io_chosenOH               (cmdArbiter_io_chosenOH[3:0]            ), //o
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  always @(*) begin
    case(readRspIndex)
      2'b00 : _zz_io_output_r_ready = io_inputs_0_r_ready;
      2'b01 : _zz_io_output_r_ready = io_inputs_1_r_ready;
      2'b10 : _zz_io_output_r_ready = io_inputs_2_r_ready;
      default : _zz_io_output_r_ready = io_inputs_3_r_ready;
    endcase
  end

  assign io_inputs_0_ar_ready = cmdArbiter_io_inputs_0_ready;
  assign io_inputs_1_ar_ready = cmdArbiter_io_inputs_1_ready;
  assign io_inputs_2_ar_ready = cmdArbiter_io_inputs_2_ready;
  assign io_inputs_3_ar_ready = cmdArbiter_io_inputs_3_ready;
  assign io_output_ar_valid = cmdArbiter_io_output_valid;
  assign io_output_ar_payload_addr = cmdArbiter_io_output_payload_addr;
  assign io_output_ar_payload_len = cmdArbiter_io_output_payload_len;
  assign io_output_ar_payload_size = cmdArbiter_io_output_payload_size;
  assign io_output_ar_payload_burst = cmdArbiter_io_output_payload_burst;
  assign io_output_ar_payload_id = {cmdArbiter_io_chosen,cmdArbiter_io_output_payload_id};
  assign readRspIndex = io_output_r_payload_id[6 : 5];
  assign readRspSels_0 = (readRspIndex == 2'b00);
  assign readRspSels_1 = (readRspIndex == 2'b01);
  assign readRspSels_2 = (readRspIndex == 2'b10);
  assign readRspSels_3 = (readRspIndex == 2'b11);
  assign io_inputs_0_r_valid = (io_output_r_valid && readRspSels_0);
  assign io_inputs_0_r_payload_data = io_output_r_payload_data;
  assign io_inputs_0_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_0_r_payload_last = io_output_r_payload_last;
  assign io_inputs_0_r_payload_id = io_output_r_payload_id[4 : 0];
  assign io_inputs_1_r_valid = (io_output_r_valid && readRspSels_1);
  assign io_inputs_1_r_payload_data = io_output_r_payload_data;
  assign io_inputs_1_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_1_r_payload_last = io_output_r_payload_last;
  assign io_inputs_1_r_payload_id = io_output_r_payload_id[4 : 0];
  assign io_inputs_2_r_valid = (io_output_r_valid && readRspSels_2);
  assign io_inputs_2_r_payload_data = io_output_r_payload_data;
  assign io_inputs_2_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_2_r_payload_last = io_output_r_payload_last;
  assign io_inputs_2_r_payload_id = io_output_r_payload_id[4 : 0];
  assign io_inputs_3_r_valid = (io_output_r_valid && readRspSels_3);
  assign io_inputs_3_r_payload_data = io_output_r_payload_data;
  assign io_inputs_3_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_3_r_payload_last = io_output_r_payload_last;
  assign io_inputs_3_r_payload_id = io_output_r_payload_id[4 : 0];
  assign io_output_r_ready = _zz_io_output_r_ready;

endmodule

//Axi4WriteOnlyDecoder_3 replaced by Axi4WriteOnlyDecoder

//Axi4ReadOnlyDecoder_3 replaced by Axi4ReadOnlyDecoder

module Axi4WriteOnlyDecoder_2 (
  input  wire          io_input_aw_valid,
  output wire          io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [2:0]    io_input_aw_payload_id,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire [2:0]    io_input_aw_payload_prot,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [31:0]   io_input_w_payload_data,
  input  wire [3:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output reg  [2:0]    io_input_b_payload_id,
  output reg  [1:0]    io_input_b_payload_resp,
  output wire          io_outputs_0_aw_valid,
  input  wire          io_outputs_0_aw_ready,
  output wire [31:0]   io_outputs_0_aw_payload_addr,
  output wire [2:0]    io_outputs_0_aw_payload_id,
  output wire [7:0]    io_outputs_0_aw_payload_len,
  output wire [2:0]    io_outputs_0_aw_payload_size,
  output wire [1:0]    io_outputs_0_aw_payload_burst,
  output wire [2:0]    io_outputs_0_aw_payload_prot,
  output wire          io_outputs_0_w_valid,
  input  wire          io_outputs_0_w_ready,
  output wire [31:0]   io_outputs_0_w_payload_data,
  output wire [3:0]    io_outputs_0_w_payload_strb,
  output wire          io_outputs_0_w_payload_last,
  input  wire          io_outputs_0_b_valid,
  output wire          io_outputs_0_b_ready,
  input  wire [2:0]    io_outputs_0_b_payload_id,
  input  wire [1:0]    io_outputs_0_b_payload_resp,
  output wire          io_outputs_1_aw_valid,
  input  wire          io_outputs_1_aw_ready,
  output wire [31:0]   io_outputs_1_aw_payload_addr,
  output wire [2:0]    io_outputs_1_aw_payload_id,
  output wire [7:0]    io_outputs_1_aw_payload_len,
  output wire [2:0]    io_outputs_1_aw_payload_size,
  output wire [1:0]    io_outputs_1_aw_payload_burst,
  output wire [2:0]    io_outputs_1_aw_payload_prot,
  output wire          io_outputs_1_w_valid,
  input  wire          io_outputs_1_w_ready,
  output wire [31:0]   io_outputs_1_w_payload_data,
  output wire [3:0]    io_outputs_1_w_payload_strb,
  output wire          io_outputs_1_w_payload_last,
  input  wire          io_outputs_1_b_valid,
  output wire          io_outputs_1_b_ready,
  input  wire [2:0]    io_outputs_1_b_payload_id,
  input  wire [1:0]    io_outputs_1_b_payload_resp,
  output wire          io_outputs_2_aw_valid,
  input  wire          io_outputs_2_aw_ready,
  output wire [31:0]   io_outputs_2_aw_payload_addr,
  output wire [2:0]    io_outputs_2_aw_payload_id,
  output wire [7:0]    io_outputs_2_aw_payload_len,
  output wire [2:0]    io_outputs_2_aw_payload_size,
  output wire [1:0]    io_outputs_2_aw_payload_burst,
  output wire [2:0]    io_outputs_2_aw_payload_prot,
  output wire          io_outputs_2_w_valid,
  input  wire          io_outputs_2_w_ready,
  output wire [31:0]   io_outputs_2_w_payload_data,
  output wire [3:0]    io_outputs_2_w_payload_strb,
  output wire          io_outputs_2_w_payload_last,
  input  wire          io_outputs_2_b_valid,
  output wire          io_outputs_2_b_ready,
  input  wire [2:0]    io_outputs_2_b_payload_id,
  input  wire [1:0]    io_outputs_2_b_payload_resp,
  input  wire          clk,
  input  wire          reset
);

  wire                errorSlave_io_axi_aw_valid;
  wire                errorSlave_io_axi_w_valid;
  wire                errorSlave_io_axi_aw_ready;
  wire                errorSlave_io_axi_w_ready;
  wire                errorSlave_io_axi_b_valid;
  wire       [2:0]    errorSlave_io_axi_b_payload_id;
  wire       [1:0]    errorSlave_io_axi_b_payload_resp;
  reg        [2:0]    _zz_io_input_b_payload_id;
  reg        [1:0]    _zz_io_input_b_payload_resp;
  wire                cmdAllowedStart;
  wire                io_input_aw_fire;
  wire                io_input_b_fire;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_mayOverflow;
  wire                pendingCmdCounter_mayUnderflow;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  wire                pendingCmdCounter_willUnderflowIfDec;
  wire                pendingCmdCounter_willUnderflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l767;
  wire                when_Utils_l769;
  wire                io_input_w_fire;
  wire                when_Utils_l735;
  reg                 pendingDataCounter_incrementIt;
  reg                 pendingDataCounter_decrementIt;
  wire       [2:0]    pendingDataCounter_valueNext;
  reg        [2:0]    pendingDataCounter_value;
  wire                pendingDataCounter_mayOverflow;
  wire                pendingDataCounter_mayUnderflow;
  wire                pendingDataCounter_willOverflowIfInc;
  wire                pendingDataCounter_willOverflow;
  wire                pendingDataCounter_willUnderflowIfDec;
  wire                pendingDataCounter_willUnderflow;
  reg        [2:0]    pendingDataCounter_finalIncrement;
  wire                when_Utils_l767_1;
  wire                when_Utils_l769_1;
  wire       [2:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [2:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                allowData;
  reg                 _zz_cmdAllowedStart;
  wire                _zz_io_outputs_1_w_valid;
  wire                _zz_io_outputs_2_w_valid;
  wire       [1:0]    writeRspIndex;

  Axi4WriteOnlyErrorSlave_2 errorSlave (
    .io_axi_aw_valid         (errorSlave_io_axi_aw_valid           ), //i
    .io_axi_aw_ready         (errorSlave_io_axi_aw_ready           ), //o
    .io_axi_aw_payload_addr  (io_input_aw_payload_addr[31:0]       ), //i
    .io_axi_aw_payload_id    (io_input_aw_payload_id[2:0]          ), //i
    .io_axi_aw_payload_len   (io_input_aw_payload_len[7:0]         ), //i
    .io_axi_aw_payload_size  (io_input_aw_payload_size[2:0]        ), //i
    .io_axi_aw_payload_burst (io_input_aw_payload_burst[1:0]       ), //i
    .io_axi_aw_payload_prot  (io_input_aw_payload_prot[2:0]        ), //i
    .io_axi_w_valid          (errorSlave_io_axi_w_valid            ), //i
    .io_axi_w_ready          (errorSlave_io_axi_w_ready            ), //o
    .io_axi_w_payload_data   (io_input_w_payload_data[31:0]        ), //i
    .io_axi_w_payload_strb   (io_input_w_payload_strb[3:0]         ), //i
    .io_axi_w_payload_last   (io_input_w_payload_last              ), //i
    .io_axi_b_valid          (errorSlave_io_axi_b_valid            ), //o
    .io_axi_b_ready          (io_input_b_ready                     ), //i
    .io_axi_b_payload_id     (errorSlave_io_axi_b_payload_id[2:0]  ), //o
    .io_axi_b_payload_resp   (errorSlave_io_axi_b_payload_resp[1:0]), //o
    .clk                     (clk                                  ), //i
    .reset                   (reset                                )  //i
  );
  always @(*) begin
    case(writeRspIndex)
      2'b00 : begin
        _zz_io_input_b_payload_id = io_outputs_0_b_payload_id;
        _zz_io_input_b_payload_resp = io_outputs_0_b_payload_resp;
      end
      2'b01 : begin
        _zz_io_input_b_payload_id = io_outputs_1_b_payload_id;
        _zz_io_input_b_payload_resp = io_outputs_1_b_payload_resp;
      end
      default : begin
        _zz_io_input_b_payload_id = io_outputs_2_b_payload_id;
        _zz_io_input_b_payload_resp = io_outputs_2_b_payload_resp;
      end
    endcase
  end

  assign io_input_aw_fire = (io_input_aw_valid && io_input_aw_ready);
  assign io_input_b_fire = (io_input_b_valid && io_input_b_ready);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_aw_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(io_input_b_fire) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_mayOverflow = (pendingCmdCounter_value == 3'b111);
  assign pendingCmdCounter_mayUnderflow = (pendingCmdCounter_value == 3'b000);
  assign pendingCmdCounter_willOverflowIfInc = (pendingCmdCounter_mayOverflow && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign pendingCmdCounter_willUnderflowIfDec = (pendingCmdCounter_mayUnderflow && (! pendingCmdCounter_incrementIt));
  assign pendingCmdCounter_willUnderflow = (pendingCmdCounter_willUnderflowIfDec && pendingCmdCounter_decrementIt);
  assign when_Utils_l767 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l767) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l769) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l769 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign io_input_w_fire = (io_input_w_valid && io_input_w_ready);
  assign when_Utils_l735 = (io_input_w_fire && io_input_w_payload_last);
  always @(*) begin
    pendingDataCounter_incrementIt = 1'b0;
    if(cmdAllowedStart) begin
      pendingDataCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingDataCounter_decrementIt = 1'b0;
    if(when_Utils_l735) begin
      pendingDataCounter_decrementIt = 1'b1;
    end
  end

  assign pendingDataCounter_mayOverflow = (pendingDataCounter_value == 3'b111);
  assign pendingDataCounter_mayUnderflow = (pendingDataCounter_value == 3'b000);
  assign pendingDataCounter_willOverflowIfInc = (pendingDataCounter_mayOverflow && (! pendingDataCounter_decrementIt));
  assign pendingDataCounter_willOverflow = (pendingDataCounter_willOverflowIfInc && pendingDataCounter_incrementIt);
  assign pendingDataCounter_willUnderflowIfDec = (pendingDataCounter_mayUnderflow && (! pendingDataCounter_incrementIt));
  assign pendingDataCounter_willUnderflow = (pendingDataCounter_willUnderflowIfDec && pendingDataCounter_decrementIt);
  assign when_Utils_l767_1 = (pendingDataCounter_incrementIt && (! pendingDataCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l767_1) begin
      pendingDataCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l769_1) begin
        pendingDataCounter_finalIncrement = 3'b111;
      end else begin
        pendingDataCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l769_1 = ((! pendingDataCounter_incrementIt) && pendingDataCounter_decrementIt);
  assign pendingDataCounter_valueNext = (pendingDataCounter_value + pendingDataCounter_finalIncrement);
  assign decodedCmdSels = {(((io_input_aw_payload_addr & (~ 32'h000003ff)) == 32'hbfd00000) && io_input_aw_valid),{(((io_input_aw_payload_addr & (~ 32'h003fffff)) == 32'h80400000) && io_input_aw_valid),(((io_input_aw_payload_addr & (~ 32'h003fffff)) == 32'h80000000) && io_input_aw_valid)}};
  assign decodedCmdError = (decodedCmdSels == 3'b000);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign allowData = (pendingDataCounter_value != 3'b000);
  assign cmdAllowedStart = ((io_input_aw_valid && allowCmd) && _zz_cmdAllowedStart);
  assign io_input_aw_ready = (((|(decodedCmdSels & {io_outputs_2_aw_ready,{io_outputs_1_aw_ready,io_outputs_0_aw_ready}})) || (decodedCmdError && errorSlave_io_axi_aw_ready)) && allowCmd);
  assign errorSlave_io_axi_aw_valid = ((io_input_aw_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_aw_valid = ((io_input_aw_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_0_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_0_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_0_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_0_aw_payload_burst = io_input_aw_payload_burst;
  assign io_outputs_0_aw_payload_prot = io_input_aw_payload_prot;
  assign io_outputs_1_aw_valid = ((io_input_aw_valid && decodedCmdSels[1]) && allowCmd);
  assign io_outputs_1_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_1_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_1_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_1_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_1_aw_payload_burst = io_input_aw_payload_burst;
  assign io_outputs_1_aw_payload_prot = io_input_aw_payload_prot;
  assign io_outputs_2_aw_valid = ((io_input_aw_valid && decodedCmdSels[2]) && allowCmd);
  assign io_outputs_2_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_2_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_2_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_2_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_2_aw_payload_burst = io_input_aw_payload_burst;
  assign io_outputs_2_aw_payload_prot = io_input_aw_payload_prot;
  assign io_input_w_ready = (((|(pendingSels & {io_outputs_2_w_ready,{io_outputs_1_w_ready,io_outputs_0_w_ready}})) || (pendingError && errorSlave_io_axi_w_ready)) && allowData);
  assign errorSlave_io_axi_w_valid = ((io_input_w_valid && pendingError) && allowData);
  assign _zz_io_outputs_1_w_valid = pendingSels[1];
  assign _zz_io_outputs_2_w_valid = pendingSels[2];
  assign io_outputs_0_w_valid = ((io_input_w_valid && pendingSels[0]) && allowData);
  assign io_outputs_0_w_payload_data = io_input_w_payload_data;
  assign io_outputs_0_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_0_w_payload_last = io_input_w_payload_last;
  assign io_outputs_1_w_valid = ((io_input_w_valid && _zz_io_outputs_1_w_valid) && allowData);
  assign io_outputs_1_w_payload_data = io_input_w_payload_data;
  assign io_outputs_1_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_1_w_payload_last = io_input_w_payload_last;
  assign io_outputs_2_w_valid = ((io_input_w_valid && _zz_io_outputs_2_w_valid) && allowData);
  assign io_outputs_2_w_payload_data = io_input_w_payload_data;
  assign io_outputs_2_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_2_w_payload_last = io_input_w_payload_last;
  assign writeRspIndex = {_zz_io_outputs_2_w_valid,_zz_io_outputs_1_w_valid};
  assign io_input_b_valid = ((|{io_outputs_2_b_valid,{io_outputs_1_b_valid,io_outputs_0_b_valid}}) || errorSlave_io_axi_b_valid);
  always @(*) begin
    io_input_b_payload_id = _zz_io_input_b_payload_id;
    if(pendingError) begin
      io_input_b_payload_id = errorSlave_io_axi_b_payload_id;
    end
  end

  always @(*) begin
    io_input_b_payload_resp = _zz_io_input_b_payload_resp;
    if(pendingError) begin
      io_input_b_payload_resp = errorSlave_io_axi_b_payload_resp;
    end
  end

  assign io_outputs_0_b_ready = io_input_b_ready;
  assign io_outputs_1_b_ready = io_input_b_ready;
  assign io_outputs_2_b_ready = io_input_b_ready;
  always @(posedge clk) begin
    if(reset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingDataCounter_value <= 3'b000;
      pendingSels <= 3'b000;
      pendingError <= 1'b0;
      _zz_cmdAllowedStart <= 1'b1;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      pendingDataCounter_value <= pendingDataCounter_valueNext;
      if(cmdAllowedStart) begin
        pendingSels <= decodedCmdSels;
      end
      if(cmdAllowedStart) begin
        pendingError <= decodedCmdError;
      end
      if(cmdAllowedStart) begin
        _zz_cmdAllowedStart <= 1'b0;
      end
      if(io_input_aw_ready) begin
        _zz_cmdAllowedStart <= 1'b1;
      end
    end
  end


endmodule

module Axi4ReadOnlyDecoder_2 (
  input  wire          io_input_ar_valid,
  output wire          io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [2:0]    io_input_ar_payload_id,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  input  wire [2:0]    io_input_ar_payload_prot,
  output reg           io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [31:0]   io_input_r_payload_data,
  output reg  [2:0]    io_input_r_payload_id,
  output reg  [1:0]    io_input_r_payload_resp,
  output reg           io_input_r_payload_last,
  output wire          io_outputs_0_ar_valid,
  input  wire          io_outputs_0_ar_ready,
  output wire [31:0]   io_outputs_0_ar_payload_addr,
  output wire [2:0]    io_outputs_0_ar_payload_id,
  output wire [7:0]    io_outputs_0_ar_payload_len,
  output wire [2:0]    io_outputs_0_ar_payload_size,
  output wire [1:0]    io_outputs_0_ar_payload_burst,
  output wire [2:0]    io_outputs_0_ar_payload_prot,
  input  wire          io_outputs_0_r_valid,
  output wire          io_outputs_0_r_ready,
  input  wire [31:0]   io_outputs_0_r_payload_data,
  input  wire [2:0]    io_outputs_0_r_payload_id,
  input  wire [1:0]    io_outputs_0_r_payload_resp,
  input  wire          io_outputs_0_r_payload_last,
  output wire          io_outputs_1_ar_valid,
  input  wire          io_outputs_1_ar_ready,
  output wire [31:0]   io_outputs_1_ar_payload_addr,
  output wire [2:0]    io_outputs_1_ar_payload_id,
  output wire [7:0]    io_outputs_1_ar_payload_len,
  output wire [2:0]    io_outputs_1_ar_payload_size,
  output wire [1:0]    io_outputs_1_ar_payload_burst,
  output wire [2:0]    io_outputs_1_ar_payload_prot,
  input  wire          io_outputs_1_r_valid,
  output wire          io_outputs_1_r_ready,
  input  wire [31:0]   io_outputs_1_r_payload_data,
  input  wire [2:0]    io_outputs_1_r_payload_id,
  input  wire [1:0]    io_outputs_1_r_payload_resp,
  input  wire          io_outputs_1_r_payload_last,
  output wire          io_outputs_2_ar_valid,
  input  wire          io_outputs_2_ar_ready,
  output wire [31:0]   io_outputs_2_ar_payload_addr,
  output wire [2:0]    io_outputs_2_ar_payload_id,
  output wire [7:0]    io_outputs_2_ar_payload_len,
  output wire [2:0]    io_outputs_2_ar_payload_size,
  output wire [1:0]    io_outputs_2_ar_payload_burst,
  output wire [2:0]    io_outputs_2_ar_payload_prot,
  input  wire          io_outputs_2_r_valid,
  output wire          io_outputs_2_r_ready,
  input  wire [31:0]   io_outputs_2_r_payload_data,
  input  wire [2:0]    io_outputs_2_r_payload_id,
  input  wire [1:0]    io_outputs_2_r_payload_resp,
  input  wire          io_outputs_2_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  wire                errorSlave_io_axi_ar_valid;
  wire                errorSlave_io_axi_ar_ready;
  wire                errorSlave_io_axi_r_valid;
  wire       [31:0]   errorSlave_io_axi_r_payload_data;
  wire       [2:0]    errorSlave_io_axi_r_payload_id;
  wire       [1:0]    errorSlave_io_axi_r_payload_resp;
  wire                errorSlave_io_axi_r_payload_last;
  reg        [31:0]   _zz_io_input_r_payload_data;
  reg        [2:0]    _zz_io_input_r_payload_id;
  reg        [1:0]    _zz_io_input_r_payload_resp;
  reg                 _zz_io_input_r_payload_last;
  wire                io_input_ar_fire;
  wire                io_input_r_fire;
  wire                when_Utils_l735;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_mayOverflow;
  wire                pendingCmdCounter_mayUnderflow;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  wire                pendingCmdCounter_willUnderflowIfDec;
  wire                pendingCmdCounter_willUnderflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l767;
  wire                when_Utils_l769;
  wire       [2:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [2:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                _zz_readRspIndex;
  wire                _zz_readRspIndex_1;
  wire       [1:0]    readRspIndex;

  Axi4ReadOnlyErrorSlave_2 errorSlave (
    .io_axi_ar_valid         (errorSlave_io_axi_ar_valid            ), //i
    .io_axi_ar_ready         (errorSlave_io_axi_ar_ready            ), //o
    .io_axi_ar_payload_addr  (io_input_ar_payload_addr[31:0]        ), //i
    .io_axi_ar_payload_id    (io_input_ar_payload_id[2:0]           ), //i
    .io_axi_ar_payload_len   (io_input_ar_payload_len[7:0]          ), //i
    .io_axi_ar_payload_size  (io_input_ar_payload_size[2:0]         ), //i
    .io_axi_ar_payload_burst (io_input_ar_payload_burst[1:0]        ), //i
    .io_axi_ar_payload_prot  (io_input_ar_payload_prot[2:0]         ), //i
    .io_axi_r_valid          (errorSlave_io_axi_r_valid             ), //o
    .io_axi_r_ready          (io_input_r_ready                      ), //i
    .io_axi_r_payload_data   (errorSlave_io_axi_r_payload_data[31:0]), //o
    .io_axi_r_payload_id     (errorSlave_io_axi_r_payload_id[2:0]   ), //o
    .io_axi_r_payload_resp   (errorSlave_io_axi_r_payload_resp[1:0] ), //o
    .io_axi_r_payload_last   (errorSlave_io_axi_r_payload_last      ), //o
    .clk                     (clk                                   ), //i
    .reset                   (reset                                 )  //i
  );
  always @(*) begin
    case(readRspIndex)
      2'b00 : begin
        _zz_io_input_r_payload_data = io_outputs_0_r_payload_data;
        _zz_io_input_r_payload_id = io_outputs_0_r_payload_id;
        _zz_io_input_r_payload_resp = io_outputs_0_r_payload_resp;
        _zz_io_input_r_payload_last = io_outputs_0_r_payload_last;
      end
      2'b01 : begin
        _zz_io_input_r_payload_data = io_outputs_1_r_payload_data;
        _zz_io_input_r_payload_id = io_outputs_1_r_payload_id;
        _zz_io_input_r_payload_resp = io_outputs_1_r_payload_resp;
        _zz_io_input_r_payload_last = io_outputs_1_r_payload_last;
      end
      default : begin
        _zz_io_input_r_payload_data = io_outputs_2_r_payload_data;
        _zz_io_input_r_payload_id = io_outputs_2_r_payload_id;
        _zz_io_input_r_payload_resp = io_outputs_2_r_payload_resp;
        _zz_io_input_r_payload_last = io_outputs_2_r_payload_last;
      end
    endcase
  end

  assign io_input_ar_fire = (io_input_ar_valid && io_input_ar_ready);
  assign io_input_r_fire = (io_input_r_valid && io_input_r_ready);
  assign when_Utils_l735 = (io_input_r_fire && io_input_r_payload_last);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_ar_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(when_Utils_l735) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_mayOverflow = (pendingCmdCounter_value == 3'b111);
  assign pendingCmdCounter_mayUnderflow = (pendingCmdCounter_value == 3'b000);
  assign pendingCmdCounter_willOverflowIfInc = (pendingCmdCounter_mayOverflow && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign pendingCmdCounter_willUnderflowIfDec = (pendingCmdCounter_mayUnderflow && (! pendingCmdCounter_incrementIt));
  assign pendingCmdCounter_willUnderflow = (pendingCmdCounter_willUnderflowIfDec && pendingCmdCounter_decrementIt);
  assign when_Utils_l767 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l767) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l769) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l769 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign decodedCmdSels = {(((io_input_ar_payload_addr & (~ 32'h000003ff)) == 32'hbfd00000) && io_input_ar_valid),{(((io_input_ar_payload_addr & (~ 32'h003fffff)) == 32'h80400000) && io_input_ar_valid),(((io_input_ar_payload_addr & (~ 32'h003fffff)) == 32'h80000000) && io_input_ar_valid)}};
  assign decodedCmdError = (decodedCmdSels == 3'b000);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign io_input_ar_ready = (((|(decodedCmdSels & {io_outputs_2_ar_ready,{io_outputs_1_ar_ready,io_outputs_0_ar_ready}})) || (decodedCmdError && errorSlave_io_axi_ar_ready)) && allowCmd);
  assign errorSlave_io_axi_ar_valid = ((io_input_ar_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_ar_valid = ((io_input_ar_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_0_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_0_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_0_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_0_ar_payload_burst = io_input_ar_payload_burst;
  assign io_outputs_0_ar_payload_prot = io_input_ar_payload_prot;
  assign io_outputs_1_ar_valid = ((io_input_ar_valid && decodedCmdSels[1]) && allowCmd);
  assign io_outputs_1_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_1_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_1_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_1_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_1_ar_payload_burst = io_input_ar_payload_burst;
  assign io_outputs_1_ar_payload_prot = io_input_ar_payload_prot;
  assign io_outputs_2_ar_valid = ((io_input_ar_valid && decodedCmdSels[2]) && allowCmd);
  assign io_outputs_2_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_2_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_2_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_2_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_2_ar_payload_burst = io_input_ar_payload_burst;
  assign io_outputs_2_ar_payload_prot = io_input_ar_payload_prot;
  assign _zz_readRspIndex = pendingSels[1];
  assign _zz_readRspIndex_1 = pendingSels[2];
  assign readRspIndex = {_zz_readRspIndex_1,_zz_readRspIndex};
  always @(*) begin
    io_input_r_valid = (|{io_outputs_2_r_valid,{io_outputs_1_r_valid,io_outputs_0_r_valid}});
    if(errorSlave_io_axi_r_valid) begin
      io_input_r_valid = 1'b1;
    end
  end

  assign io_input_r_payload_data = _zz_io_input_r_payload_data;
  always @(*) begin
    io_input_r_payload_id = _zz_io_input_r_payload_id;
    if(pendingError) begin
      io_input_r_payload_id = errorSlave_io_axi_r_payload_id;
    end
  end

  always @(*) begin
    io_input_r_payload_resp = _zz_io_input_r_payload_resp;
    if(pendingError) begin
      io_input_r_payload_resp = errorSlave_io_axi_r_payload_resp;
    end
  end

  always @(*) begin
    io_input_r_payload_last = _zz_io_input_r_payload_last;
    if(pendingError) begin
      io_input_r_payload_last = errorSlave_io_axi_r_payload_last;
    end
  end

  assign io_outputs_0_r_ready = io_input_r_ready;
  assign io_outputs_1_r_ready = io_input_r_ready;
  assign io_outputs_2_r_ready = io_input_r_ready;
  always @(posedge clk) begin
    if(reset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingSels <= 3'b000;
      pendingError <= 1'b0;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      if(io_input_ar_ready) begin
        pendingSels <= decodedCmdSels;
      end
      if(io_input_ar_ready) begin
        pendingError <= decodedCmdError;
      end
    end
  end


endmodule

//Axi4WriteOnlyDecoder_1 replaced by Axi4WriteOnlyDecoder

//Axi4ReadOnlyDecoder_1 replaced by Axi4ReadOnlyDecoder

module Axi4WriteOnlyDecoder (
  input  wire          io_input_aw_valid,
  output wire          io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [3:0]    io_input_aw_payload_id,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [31:0]   io_input_w_payload_data,
  input  wire [3:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output reg  [3:0]    io_input_b_payload_id,
  output reg  [1:0]    io_input_b_payload_resp,
  output wire          io_outputs_0_aw_valid,
  input  wire          io_outputs_0_aw_ready,
  output wire [31:0]   io_outputs_0_aw_payload_addr,
  output wire [3:0]    io_outputs_0_aw_payload_id,
  output wire [7:0]    io_outputs_0_aw_payload_len,
  output wire [2:0]    io_outputs_0_aw_payload_size,
  output wire [1:0]    io_outputs_0_aw_payload_burst,
  output wire          io_outputs_0_w_valid,
  input  wire          io_outputs_0_w_ready,
  output wire [31:0]   io_outputs_0_w_payload_data,
  output wire [3:0]    io_outputs_0_w_payload_strb,
  output wire          io_outputs_0_w_payload_last,
  input  wire          io_outputs_0_b_valid,
  output wire          io_outputs_0_b_ready,
  input  wire [3:0]    io_outputs_0_b_payload_id,
  input  wire [1:0]    io_outputs_0_b_payload_resp,
  output wire          io_outputs_1_aw_valid,
  input  wire          io_outputs_1_aw_ready,
  output wire [31:0]   io_outputs_1_aw_payload_addr,
  output wire [3:0]    io_outputs_1_aw_payload_id,
  output wire [7:0]    io_outputs_1_aw_payload_len,
  output wire [2:0]    io_outputs_1_aw_payload_size,
  output wire [1:0]    io_outputs_1_aw_payload_burst,
  output wire          io_outputs_1_w_valid,
  input  wire          io_outputs_1_w_ready,
  output wire [31:0]   io_outputs_1_w_payload_data,
  output wire [3:0]    io_outputs_1_w_payload_strb,
  output wire          io_outputs_1_w_payload_last,
  input  wire          io_outputs_1_b_valid,
  output wire          io_outputs_1_b_ready,
  input  wire [3:0]    io_outputs_1_b_payload_id,
  input  wire [1:0]    io_outputs_1_b_payload_resp,
  output wire          io_outputs_2_aw_valid,
  input  wire          io_outputs_2_aw_ready,
  output wire [31:0]   io_outputs_2_aw_payload_addr,
  output wire [3:0]    io_outputs_2_aw_payload_id,
  output wire [7:0]    io_outputs_2_aw_payload_len,
  output wire [2:0]    io_outputs_2_aw_payload_size,
  output wire [1:0]    io_outputs_2_aw_payload_burst,
  output wire          io_outputs_2_w_valid,
  input  wire          io_outputs_2_w_ready,
  output wire [31:0]   io_outputs_2_w_payload_data,
  output wire [3:0]    io_outputs_2_w_payload_strb,
  output wire          io_outputs_2_w_payload_last,
  input  wire          io_outputs_2_b_valid,
  output wire          io_outputs_2_b_ready,
  input  wire [3:0]    io_outputs_2_b_payload_id,
  input  wire [1:0]    io_outputs_2_b_payload_resp,
  input  wire          clk,
  input  wire          reset
);

  wire                errorSlave_io_axi_aw_valid;
  wire                errorSlave_io_axi_w_valid;
  wire                errorSlave_io_axi_aw_ready;
  wire                errorSlave_io_axi_w_ready;
  wire                errorSlave_io_axi_b_valid;
  wire       [3:0]    errorSlave_io_axi_b_payload_id;
  wire       [1:0]    errorSlave_io_axi_b_payload_resp;
  reg        [3:0]    _zz_io_input_b_payload_id;
  reg        [1:0]    _zz_io_input_b_payload_resp;
  wire                cmdAllowedStart;
  wire                io_input_aw_fire;
  wire                io_input_b_fire;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_mayOverflow;
  wire                pendingCmdCounter_mayUnderflow;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  wire                pendingCmdCounter_willUnderflowIfDec;
  wire                pendingCmdCounter_willUnderflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l767;
  wire                when_Utils_l769;
  wire                io_input_w_fire;
  wire                when_Utils_l735;
  reg                 pendingDataCounter_incrementIt;
  reg                 pendingDataCounter_decrementIt;
  wire       [2:0]    pendingDataCounter_valueNext;
  reg        [2:0]    pendingDataCounter_value;
  wire                pendingDataCounter_mayOverflow;
  wire                pendingDataCounter_mayUnderflow;
  wire                pendingDataCounter_willOverflowIfInc;
  wire                pendingDataCounter_willOverflow;
  wire                pendingDataCounter_willUnderflowIfDec;
  wire                pendingDataCounter_willUnderflow;
  reg        [2:0]    pendingDataCounter_finalIncrement;
  wire                when_Utils_l767_1;
  wire                when_Utils_l769_1;
  wire       [2:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [2:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                allowData;
  reg                 _zz_cmdAllowedStart;
  wire                _zz_io_outputs_1_w_valid;
  wire                _zz_io_outputs_2_w_valid;
  wire       [1:0]    writeRspIndex;

  Axi4WriteOnlyErrorSlave errorSlave (
    .io_axi_aw_valid         (errorSlave_io_axi_aw_valid           ), //i
    .io_axi_aw_ready         (errorSlave_io_axi_aw_ready           ), //o
    .io_axi_aw_payload_addr  (io_input_aw_payload_addr[31:0]       ), //i
    .io_axi_aw_payload_id    (io_input_aw_payload_id[3:0]          ), //i
    .io_axi_aw_payload_len   (io_input_aw_payload_len[7:0]         ), //i
    .io_axi_aw_payload_size  (io_input_aw_payload_size[2:0]        ), //i
    .io_axi_aw_payload_burst (io_input_aw_payload_burst[1:0]       ), //i
    .io_axi_w_valid          (errorSlave_io_axi_w_valid            ), //i
    .io_axi_w_ready          (errorSlave_io_axi_w_ready            ), //o
    .io_axi_w_payload_data   (io_input_w_payload_data[31:0]        ), //i
    .io_axi_w_payload_strb   (io_input_w_payload_strb[3:0]         ), //i
    .io_axi_w_payload_last   (io_input_w_payload_last              ), //i
    .io_axi_b_valid          (errorSlave_io_axi_b_valid            ), //o
    .io_axi_b_ready          (io_input_b_ready                     ), //i
    .io_axi_b_payload_id     (errorSlave_io_axi_b_payload_id[3:0]  ), //o
    .io_axi_b_payload_resp   (errorSlave_io_axi_b_payload_resp[1:0]), //o
    .clk                     (clk                                  ), //i
    .reset                   (reset                                )  //i
  );
  always @(*) begin
    case(writeRspIndex)
      2'b00 : begin
        _zz_io_input_b_payload_id = io_outputs_0_b_payload_id;
        _zz_io_input_b_payload_resp = io_outputs_0_b_payload_resp;
      end
      2'b01 : begin
        _zz_io_input_b_payload_id = io_outputs_1_b_payload_id;
        _zz_io_input_b_payload_resp = io_outputs_1_b_payload_resp;
      end
      default : begin
        _zz_io_input_b_payload_id = io_outputs_2_b_payload_id;
        _zz_io_input_b_payload_resp = io_outputs_2_b_payload_resp;
      end
    endcase
  end

  assign io_input_aw_fire = (io_input_aw_valid && io_input_aw_ready);
  assign io_input_b_fire = (io_input_b_valid && io_input_b_ready);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_aw_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(io_input_b_fire) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_mayOverflow = (pendingCmdCounter_value == 3'b111);
  assign pendingCmdCounter_mayUnderflow = (pendingCmdCounter_value == 3'b000);
  assign pendingCmdCounter_willOverflowIfInc = (pendingCmdCounter_mayOverflow && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign pendingCmdCounter_willUnderflowIfDec = (pendingCmdCounter_mayUnderflow && (! pendingCmdCounter_incrementIt));
  assign pendingCmdCounter_willUnderflow = (pendingCmdCounter_willUnderflowIfDec && pendingCmdCounter_decrementIt);
  assign when_Utils_l767 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l767) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l769) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l769 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign io_input_w_fire = (io_input_w_valid && io_input_w_ready);
  assign when_Utils_l735 = (io_input_w_fire && io_input_w_payload_last);
  always @(*) begin
    pendingDataCounter_incrementIt = 1'b0;
    if(cmdAllowedStart) begin
      pendingDataCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingDataCounter_decrementIt = 1'b0;
    if(when_Utils_l735) begin
      pendingDataCounter_decrementIt = 1'b1;
    end
  end

  assign pendingDataCounter_mayOverflow = (pendingDataCounter_value == 3'b111);
  assign pendingDataCounter_mayUnderflow = (pendingDataCounter_value == 3'b000);
  assign pendingDataCounter_willOverflowIfInc = (pendingDataCounter_mayOverflow && (! pendingDataCounter_decrementIt));
  assign pendingDataCounter_willOverflow = (pendingDataCounter_willOverflowIfInc && pendingDataCounter_incrementIt);
  assign pendingDataCounter_willUnderflowIfDec = (pendingDataCounter_mayUnderflow && (! pendingDataCounter_incrementIt));
  assign pendingDataCounter_willUnderflow = (pendingDataCounter_willUnderflowIfDec && pendingDataCounter_decrementIt);
  assign when_Utils_l767_1 = (pendingDataCounter_incrementIt && (! pendingDataCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l767_1) begin
      pendingDataCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l769_1) begin
        pendingDataCounter_finalIncrement = 3'b111;
      end else begin
        pendingDataCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l769_1 = ((! pendingDataCounter_incrementIt) && pendingDataCounter_decrementIt);
  assign pendingDataCounter_valueNext = (pendingDataCounter_value + pendingDataCounter_finalIncrement);
  assign decodedCmdSels = {(((io_input_aw_payload_addr & (~ 32'h000003ff)) == 32'hbfd00000) && io_input_aw_valid),{(((io_input_aw_payload_addr & (~ 32'h003fffff)) == 32'h80400000) && io_input_aw_valid),(((io_input_aw_payload_addr & (~ 32'h003fffff)) == 32'h80000000) && io_input_aw_valid)}};
  assign decodedCmdError = (decodedCmdSels == 3'b000);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign allowData = (pendingDataCounter_value != 3'b000);
  assign cmdAllowedStart = ((io_input_aw_valid && allowCmd) && _zz_cmdAllowedStart);
  assign io_input_aw_ready = (((|(decodedCmdSels & {io_outputs_2_aw_ready,{io_outputs_1_aw_ready,io_outputs_0_aw_ready}})) || (decodedCmdError && errorSlave_io_axi_aw_ready)) && allowCmd);
  assign errorSlave_io_axi_aw_valid = ((io_input_aw_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_aw_valid = ((io_input_aw_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_0_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_0_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_0_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_0_aw_payload_burst = io_input_aw_payload_burst;
  assign io_outputs_1_aw_valid = ((io_input_aw_valid && decodedCmdSels[1]) && allowCmd);
  assign io_outputs_1_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_1_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_1_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_1_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_1_aw_payload_burst = io_input_aw_payload_burst;
  assign io_outputs_2_aw_valid = ((io_input_aw_valid && decodedCmdSels[2]) && allowCmd);
  assign io_outputs_2_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_2_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_2_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_2_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_2_aw_payload_burst = io_input_aw_payload_burst;
  assign io_input_w_ready = (((|(pendingSels & {io_outputs_2_w_ready,{io_outputs_1_w_ready,io_outputs_0_w_ready}})) || (pendingError && errorSlave_io_axi_w_ready)) && allowData);
  assign errorSlave_io_axi_w_valid = ((io_input_w_valid && pendingError) && allowData);
  assign _zz_io_outputs_1_w_valid = pendingSels[1];
  assign _zz_io_outputs_2_w_valid = pendingSels[2];
  assign io_outputs_0_w_valid = ((io_input_w_valid && pendingSels[0]) && allowData);
  assign io_outputs_0_w_payload_data = io_input_w_payload_data;
  assign io_outputs_0_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_0_w_payload_last = io_input_w_payload_last;
  assign io_outputs_1_w_valid = ((io_input_w_valid && _zz_io_outputs_1_w_valid) && allowData);
  assign io_outputs_1_w_payload_data = io_input_w_payload_data;
  assign io_outputs_1_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_1_w_payload_last = io_input_w_payload_last;
  assign io_outputs_2_w_valid = ((io_input_w_valid && _zz_io_outputs_2_w_valid) && allowData);
  assign io_outputs_2_w_payload_data = io_input_w_payload_data;
  assign io_outputs_2_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_2_w_payload_last = io_input_w_payload_last;
  assign writeRspIndex = {_zz_io_outputs_2_w_valid,_zz_io_outputs_1_w_valid};
  assign io_input_b_valid = ((|{io_outputs_2_b_valid,{io_outputs_1_b_valid,io_outputs_0_b_valid}}) || errorSlave_io_axi_b_valid);
  always @(*) begin
    io_input_b_payload_id = _zz_io_input_b_payload_id;
    if(pendingError) begin
      io_input_b_payload_id = errorSlave_io_axi_b_payload_id;
    end
  end

  always @(*) begin
    io_input_b_payload_resp = _zz_io_input_b_payload_resp;
    if(pendingError) begin
      io_input_b_payload_resp = errorSlave_io_axi_b_payload_resp;
    end
  end

  assign io_outputs_0_b_ready = io_input_b_ready;
  assign io_outputs_1_b_ready = io_input_b_ready;
  assign io_outputs_2_b_ready = io_input_b_ready;
  always @(posedge clk) begin
    if(reset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingDataCounter_value <= 3'b000;
      pendingSels <= 3'b000;
      pendingError <= 1'b0;
      _zz_cmdAllowedStart <= 1'b1;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      pendingDataCounter_value <= pendingDataCounter_valueNext;
      if(cmdAllowedStart) begin
        pendingSels <= decodedCmdSels;
      end
      if(cmdAllowedStart) begin
        pendingError <= decodedCmdError;
      end
      if(cmdAllowedStart) begin
        _zz_cmdAllowedStart <= 1'b0;
      end
      if(io_input_aw_ready) begin
        _zz_cmdAllowedStart <= 1'b1;
      end
    end
  end


endmodule

module Axi4ReadOnlyDecoder (
  input  wire          io_input_ar_valid,
  output wire          io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [3:0]    io_input_ar_payload_id,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  output reg           io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [31:0]   io_input_r_payload_data,
  output reg  [3:0]    io_input_r_payload_id,
  output reg  [1:0]    io_input_r_payload_resp,
  output reg           io_input_r_payload_last,
  output wire          io_outputs_0_ar_valid,
  input  wire          io_outputs_0_ar_ready,
  output wire [31:0]   io_outputs_0_ar_payload_addr,
  output wire [3:0]    io_outputs_0_ar_payload_id,
  output wire [7:0]    io_outputs_0_ar_payload_len,
  output wire [2:0]    io_outputs_0_ar_payload_size,
  output wire [1:0]    io_outputs_0_ar_payload_burst,
  input  wire          io_outputs_0_r_valid,
  output wire          io_outputs_0_r_ready,
  input  wire [31:0]   io_outputs_0_r_payload_data,
  input  wire [3:0]    io_outputs_0_r_payload_id,
  input  wire [1:0]    io_outputs_0_r_payload_resp,
  input  wire          io_outputs_0_r_payload_last,
  output wire          io_outputs_1_ar_valid,
  input  wire          io_outputs_1_ar_ready,
  output wire [31:0]   io_outputs_1_ar_payload_addr,
  output wire [3:0]    io_outputs_1_ar_payload_id,
  output wire [7:0]    io_outputs_1_ar_payload_len,
  output wire [2:0]    io_outputs_1_ar_payload_size,
  output wire [1:0]    io_outputs_1_ar_payload_burst,
  input  wire          io_outputs_1_r_valid,
  output wire          io_outputs_1_r_ready,
  input  wire [31:0]   io_outputs_1_r_payload_data,
  input  wire [3:0]    io_outputs_1_r_payload_id,
  input  wire [1:0]    io_outputs_1_r_payload_resp,
  input  wire          io_outputs_1_r_payload_last,
  output wire          io_outputs_2_ar_valid,
  input  wire          io_outputs_2_ar_ready,
  output wire [31:0]   io_outputs_2_ar_payload_addr,
  output wire [3:0]    io_outputs_2_ar_payload_id,
  output wire [7:0]    io_outputs_2_ar_payload_len,
  output wire [2:0]    io_outputs_2_ar_payload_size,
  output wire [1:0]    io_outputs_2_ar_payload_burst,
  input  wire          io_outputs_2_r_valid,
  output wire          io_outputs_2_r_ready,
  input  wire [31:0]   io_outputs_2_r_payload_data,
  input  wire [3:0]    io_outputs_2_r_payload_id,
  input  wire [1:0]    io_outputs_2_r_payload_resp,
  input  wire          io_outputs_2_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  wire                errorSlave_io_axi_ar_valid;
  wire                errorSlave_io_axi_ar_ready;
  wire                errorSlave_io_axi_r_valid;
  wire       [31:0]   errorSlave_io_axi_r_payload_data;
  wire       [3:0]    errorSlave_io_axi_r_payload_id;
  wire       [1:0]    errorSlave_io_axi_r_payload_resp;
  wire                errorSlave_io_axi_r_payload_last;
  reg        [31:0]   _zz_io_input_r_payload_data;
  reg        [3:0]    _zz_io_input_r_payload_id;
  reg        [1:0]    _zz_io_input_r_payload_resp;
  reg                 _zz_io_input_r_payload_last;
  wire                io_input_ar_fire;
  wire                io_input_r_fire;
  wire                when_Utils_l735;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_mayOverflow;
  wire                pendingCmdCounter_mayUnderflow;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  wire                pendingCmdCounter_willUnderflowIfDec;
  wire                pendingCmdCounter_willUnderflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l767;
  wire                when_Utils_l769;
  wire       [2:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [2:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                _zz_readRspIndex;
  wire                _zz_readRspIndex_1;
  wire       [1:0]    readRspIndex;

  Axi4ReadOnlyErrorSlave errorSlave (
    .io_axi_ar_valid         (errorSlave_io_axi_ar_valid            ), //i
    .io_axi_ar_ready         (errorSlave_io_axi_ar_ready            ), //o
    .io_axi_ar_payload_addr  (io_input_ar_payload_addr[31:0]        ), //i
    .io_axi_ar_payload_id    (io_input_ar_payload_id[3:0]           ), //i
    .io_axi_ar_payload_len   (io_input_ar_payload_len[7:0]          ), //i
    .io_axi_ar_payload_size  (io_input_ar_payload_size[2:0]         ), //i
    .io_axi_ar_payload_burst (io_input_ar_payload_burst[1:0]        ), //i
    .io_axi_r_valid          (errorSlave_io_axi_r_valid             ), //o
    .io_axi_r_ready          (io_input_r_ready                      ), //i
    .io_axi_r_payload_data   (errorSlave_io_axi_r_payload_data[31:0]), //o
    .io_axi_r_payload_id     (errorSlave_io_axi_r_payload_id[3:0]   ), //o
    .io_axi_r_payload_resp   (errorSlave_io_axi_r_payload_resp[1:0] ), //o
    .io_axi_r_payload_last   (errorSlave_io_axi_r_payload_last      ), //o
    .clk                     (clk                                   ), //i
    .reset                   (reset                                 )  //i
  );
  always @(*) begin
    case(readRspIndex)
      2'b00 : begin
        _zz_io_input_r_payload_data = io_outputs_0_r_payload_data;
        _zz_io_input_r_payload_id = io_outputs_0_r_payload_id;
        _zz_io_input_r_payload_resp = io_outputs_0_r_payload_resp;
        _zz_io_input_r_payload_last = io_outputs_0_r_payload_last;
      end
      2'b01 : begin
        _zz_io_input_r_payload_data = io_outputs_1_r_payload_data;
        _zz_io_input_r_payload_id = io_outputs_1_r_payload_id;
        _zz_io_input_r_payload_resp = io_outputs_1_r_payload_resp;
        _zz_io_input_r_payload_last = io_outputs_1_r_payload_last;
      end
      default : begin
        _zz_io_input_r_payload_data = io_outputs_2_r_payload_data;
        _zz_io_input_r_payload_id = io_outputs_2_r_payload_id;
        _zz_io_input_r_payload_resp = io_outputs_2_r_payload_resp;
        _zz_io_input_r_payload_last = io_outputs_2_r_payload_last;
      end
    endcase
  end

  assign io_input_ar_fire = (io_input_ar_valid && io_input_ar_ready);
  assign io_input_r_fire = (io_input_r_valid && io_input_r_ready);
  assign when_Utils_l735 = (io_input_r_fire && io_input_r_payload_last);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_ar_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(when_Utils_l735) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_mayOverflow = (pendingCmdCounter_value == 3'b111);
  assign pendingCmdCounter_mayUnderflow = (pendingCmdCounter_value == 3'b000);
  assign pendingCmdCounter_willOverflowIfInc = (pendingCmdCounter_mayOverflow && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign pendingCmdCounter_willUnderflowIfDec = (pendingCmdCounter_mayUnderflow && (! pendingCmdCounter_incrementIt));
  assign pendingCmdCounter_willUnderflow = (pendingCmdCounter_willUnderflowIfDec && pendingCmdCounter_decrementIt);
  assign when_Utils_l767 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l767) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l769) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l769 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign decodedCmdSels = {(((io_input_ar_payload_addr & (~ 32'h000003ff)) == 32'hbfd00000) && io_input_ar_valid),{(((io_input_ar_payload_addr & (~ 32'h003fffff)) == 32'h80400000) && io_input_ar_valid),(((io_input_ar_payload_addr & (~ 32'h003fffff)) == 32'h80000000) && io_input_ar_valid)}};
  assign decodedCmdError = (decodedCmdSels == 3'b000);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign io_input_ar_ready = (((|(decodedCmdSels & {io_outputs_2_ar_ready,{io_outputs_1_ar_ready,io_outputs_0_ar_ready}})) || (decodedCmdError && errorSlave_io_axi_ar_ready)) && allowCmd);
  assign errorSlave_io_axi_ar_valid = ((io_input_ar_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_ar_valid = ((io_input_ar_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_0_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_0_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_0_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_0_ar_payload_burst = io_input_ar_payload_burst;
  assign io_outputs_1_ar_valid = ((io_input_ar_valid && decodedCmdSels[1]) && allowCmd);
  assign io_outputs_1_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_1_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_1_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_1_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_1_ar_payload_burst = io_input_ar_payload_burst;
  assign io_outputs_2_ar_valid = ((io_input_ar_valid && decodedCmdSels[2]) && allowCmd);
  assign io_outputs_2_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_2_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_2_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_2_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_2_ar_payload_burst = io_input_ar_payload_burst;
  assign _zz_readRspIndex = pendingSels[1];
  assign _zz_readRspIndex_1 = pendingSels[2];
  assign readRspIndex = {_zz_readRspIndex_1,_zz_readRspIndex};
  always @(*) begin
    io_input_r_valid = (|{io_outputs_2_r_valid,{io_outputs_1_r_valid,io_outputs_0_r_valid}});
    if(errorSlave_io_axi_r_valid) begin
      io_input_r_valid = 1'b1;
    end
  end

  assign io_input_r_payload_data = _zz_io_input_r_payload_data;
  always @(*) begin
    io_input_r_payload_id = _zz_io_input_r_payload_id;
    if(pendingError) begin
      io_input_r_payload_id = errorSlave_io_axi_r_payload_id;
    end
  end

  always @(*) begin
    io_input_r_payload_resp = _zz_io_input_r_payload_resp;
    if(pendingError) begin
      io_input_r_payload_resp = errorSlave_io_axi_r_payload_resp;
    end
  end

  always @(*) begin
    io_input_r_payload_last = _zz_io_input_r_payload_last;
    if(pendingError) begin
      io_input_r_payload_last = errorSlave_io_axi_r_payload_last;
    end
  end

  assign io_outputs_0_r_ready = io_input_r_ready;
  assign io_outputs_1_r_ready = io_input_r_ready;
  assign io_outputs_2_r_ready = io_input_r_ready;
  always @(posedge clk) begin
    if(reset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingSels <= 3'b000;
      pendingError <= 1'b0;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      if(io_input_ar_ready) begin
        pendingSels <= decodedCmdSels;
      end
      if(io_input_ar_ready) begin
        pendingError <= decodedCmdError;
      end
    end
  end


endmodule

//SplitGmbToAxi4Bridge_1 replaced by SplitGmbToAxi4Bridge

module SplitGmbToAxi4Bridge (
  input  wire          io_gmbIn_read_cmd_valid,
  output wire          io_gmbIn_read_cmd_ready,
  input  wire [31:0]   io_gmbIn_read_cmd_payload_address,
  input  wire [3:0]    io_gmbIn_read_cmd_payload_id,
  output wire          io_gmbIn_read_rsp_valid,
  input  wire          io_gmbIn_read_rsp_ready,
  output wire [31:0]   io_gmbIn_read_rsp_payload_data,
  output wire          io_gmbIn_read_rsp_payload_error,
  output wire [3:0]    io_gmbIn_read_rsp_payload_id,
  input  wire          io_gmbIn_write_cmd_valid,
  output wire          io_gmbIn_write_cmd_ready,
  input  wire [31:0]   io_gmbIn_write_cmd_payload_address,
  input  wire [31:0]   io_gmbIn_write_cmd_payload_data,
  input  wire [3:0]    io_gmbIn_write_cmd_payload_byteEnables,
  input  wire [3:0]    io_gmbIn_write_cmd_payload_id,
  input  wire          io_gmbIn_write_cmd_payload_last,
  output wire          io_gmbIn_write_rsp_valid,
  input  wire          io_gmbIn_write_rsp_ready,
  output wire          io_gmbIn_write_rsp_payload_error,
  output wire [3:0]    io_gmbIn_write_rsp_payload_id,
  output wire          io_axiOut_aw_valid,
  input  wire          io_axiOut_aw_ready,
  output wire [31:0]   io_axiOut_aw_payload_addr,
  output wire [3:0]    io_axiOut_aw_payload_id,
  output wire [7:0]    io_axiOut_aw_payload_len,
  output wire [2:0]    io_axiOut_aw_payload_size,
  output wire [1:0]    io_axiOut_aw_payload_burst,
  output wire          io_axiOut_w_valid,
  input  wire          io_axiOut_w_ready,
  output wire [31:0]   io_axiOut_w_payload_data,
  output wire [3:0]    io_axiOut_w_payload_strb,
  output wire          io_axiOut_w_payload_last,
  input  wire          io_axiOut_b_valid,
  output wire          io_axiOut_b_ready,
  input  wire [3:0]    io_axiOut_b_payload_id,
  input  wire [1:0]    io_axiOut_b_payload_resp,
  output wire          io_axiOut_ar_valid,
  input  wire          io_axiOut_ar_ready,
  output wire [31:0]   io_axiOut_ar_payload_addr,
  output wire [3:0]    io_axiOut_ar_payload_id,
  output wire [7:0]    io_axiOut_ar_payload_len,
  output wire [2:0]    io_axiOut_ar_payload_size,
  output wire [1:0]    io_axiOut_ar_payload_burst,
  input  wire          io_axiOut_r_valid,
  output wire          io_axiOut_r_ready,
  input  wire [31:0]   io_axiOut_r_payload_data,
  input  wire [3:0]    io_axiOut_r_payload_id,
  input  wire [1:0]    io_axiOut_r_payload_resp,
  input  wire          io_axiOut_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  wire                io_gmbIn_read_cmd_fifo_io_push_ready;
  wire                io_gmbIn_read_cmd_fifo_io_pop_valid;
  wire       [31:0]   io_gmbIn_read_cmd_fifo_io_pop_payload_address;
  wire       [3:0]    io_gmbIn_read_cmd_fifo_io_pop_payload_id;
  wire       [1:0]    io_gmbIn_read_cmd_fifo_io_occupancy;
  wire       [1:0]    io_gmbIn_read_cmd_fifo_io_availability;
  wire                io_axiOut_r_fifo_io_push_ready;
  wire                io_axiOut_r_fifo_io_pop_valid;
  wire       [31:0]   io_axiOut_r_fifo_io_pop_payload_data;
  wire       [3:0]    io_axiOut_r_fifo_io_pop_payload_id;
  wire       [1:0]    io_axiOut_r_fifo_io_pop_payload_resp;
  wire                io_axiOut_r_fifo_io_pop_payload_last;
  wire       [1:0]    io_axiOut_r_fifo_io_occupancy;
  wire       [1:0]    io_axiOut_r_fifo_io_availability;
  wire                io_gmbIn_write_cmd_fifo_io_push_ready;
  wire                io_gmbIn_write_cmd_fifo_io_pop_valid;
  wire       [31:0]   io_gmbIn_write_cmd_fifo_io_pop_payload_address;
  wire       [31:0]   io_gmbIn_write_cmd_fifo_io_pop_payload_data;
  wire       [3:0]    io_gmbIn_write_cmd_fifo_io_pop_payload_byteEnables;
  wire       [3:0]    io_gmbIn_write_cmd_fifo_io_pop_payload_id;
  wire                io_gmbIn_write_cmd_fifo_io_pop_payload_last;
  wire       [1:0]    io_gmbIn_write_cmd_fifo_io_occupancy;
  wire       [1:0]    io_gmbIn_write_cmd_fifo_io_availability;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_input_ready;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_valid;
  wire       [31:0]   io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_address;
  wire       [31:0]   io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_data;
  wire       [3:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_byteEnables;
  wire       [3:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_id;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_last;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_valid;
  wire       [31:0]   io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_address;
  wire       [31:0]   io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_data;
  wire       [3:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_byteEnables;
  wire       [3:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_id;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_last;
  wire                io_axiOut_b_fifo_io_push_ready;
  wire                io_axiOut_b_fifo_io_pop_valid;
  wire       [3:0]    io_axiOut_b_fifo_io_pop_payload_id;
  wire       [1:0]    io_axiOut_b_fifo_io_pop_payload_resp;
  wire       [1:0]    io_axiOut_b_fifo_io_occupancy;
  wire       [1:0]    io_axiOut_b_fifo_io_availability;
  wire                io_gmbIn_read_cmd_fifo_io_pop_translated_valid;
  wire                io_gmbIn_read_cmd_fifo_io_pop_translated_ready;
  wire       [31:0]   io_gmbIn_read_cmd_fifo_io_pop_translated_payload_addr;
  wire       [3:0]    io_gmbIn_read_cmd_fifo_io_pop_translated_payload_id;
  wire       [7:0]    io_gmbIn_read_cmd_fifo_io_pop_translated_payload_len;
  wire       [2:0]    io_gmbIn_read_cmd_fifo_io_pop_translated_payload_size;
  wire       [1:0]    io_gmbIn_read_cmd_fifo_io_pop_translated_payload_burst;
  wire                io_axiOut_r_fifo_io_pop_translated_valid;
  wire                io_axiOut_r_fifo_io_pop_translated_ready;
  wire       [31:0]   io_axiOut_r_fifo_io_pop_translated_payload_data;
  wire                io_axiOut_r_fifo_io_pop_translated_payload_error;
  wire       [3:0]    io_axiOut_r_fifo_io_pop_translated_payload_id;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_valid;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_ready;
  wire       [31:0]   io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_addr;
  wire       [3:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_id;
  wire       [7:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_len;
  wire       [2:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_size;
  wire       [1:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_burst;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_valid;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_ready;
  wire       [31:0]   io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_data;
  wire       [3:0]    io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_strb;
  wire                io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_last;
  wire                io_axiOut_b_fifo_io_pop_translated_valid;
  wire                io_axiOut_b_fifo_io_pop_translated_ready;
  wire                io_axiOut_b_fifo_io_pop_translated_payload_error;
  wire       [3:0]    io_axiOut_b_fifo_io_pop_translated_payload_id;

  StreamFifo io_gmbIn_read_cmd_fifo (
    .io_push_valid           (io_gmbIn_read_cmd_valid                            ), //i
    .io_push_ready           (io_gmbIn_read_cmd_fifo_io_push_ready               ), //o
    .io_push_payload_address (io_gmbIn_read_cmd_payload_address[31:0]            ), //i
    .io_push_payload_id      (io_gmbIn_read_cmd_payload_id[3:0]                  ), //i
    .io_pop_valid            (io_gmbIn_read_cmd_fifo_io_pop_valid                ), //o
    .io_pop_ready            (io_gmbIn_read_cmd_fifo_io_pop_translated_ready     ), //i
    .io_pop_payload_address  (io_gmbIn_read_cmd_fifo_io_pop_payload_address[31:0]), //o
    .io_pop_payload_id       (io_gmbIn_read_cmd_fifo_io_pop_payload_id[3:0]      ), //o
    .io_flush                (1'b0                                               ), //i
    .io_occupancy            (io_gmbIn_read_cmd_fifo_io_occupancy[1:0]           ), //o
    .io_availability         (io_gmbIn_read_cmd_fifo_io_availability[1:0]        ), //o
    .clk                     (clk                                                ), //i
    .reset                   (reset                                              )  //i
  );
  StreamFifo_1 io_axiOut_r_fifo (
    .io_push_valid        (io_axiOut_r_valid                         ), //i
    .io_push_ready        (io_axiOut_r_fifo_io_push_ready            ), //o
    .io_push_payload_data (io_axiOut_r_payload_data[31:0]            ), //i
    .io_push_payload_id   (io_axiOut_r_payload_id[3:0]               ), //i
    .io_push_payload_resp (io_axiOut_r_payload_resp[1:0]             ), //i
    .io_push_payload_last (io_axiOut_r_payload_last                  ), //i
    .io_pop_valid         (io_axiOut_r_fifo_io_pop_valid             ), //o
    .io_pop_ready         (io_axiOut_r_fifo_io_pop_translated_ready  ), //i
    .io_pop_payload_data  (io_axiOut_r_fifo_io_pop_payload_data[31:0]), //o
    .io_pop_payload_id    (io_axiOut_r_fifo_io_pop_payload_id[3:0]   ), //o
    .io_pop_payload_resp  (io_axiOut_r_fifo_io_pop_payload_resp[1:0] ), //o
    .io_pop_payload_last  (io_axiOut_r_fifo_io_pop_payload_last      ), //o
    .io_flush             (1'b0                                      ), //i
    .io_occupancy         (io_axiOut_r_fifo_io_occupancy[1:0]        ), //o
    .io_availability      (io_axiOut_r_fifo_io_availability[1:0]     ), //o
    .clk                  (clk                                       ), //i
    .reset                (reset                                     )  //i
  );
  StreamFifo_2 io_gmbIn_write_cmd_fifo (
    .io_push_valid               (io_gmbIn_write_cmd_valid                               ), //i
    .io_push_ready               (io_gmbIn_write_cmd_fifo_io_push_ready                  ), //o
    .io_push_payload_address     (io_gmbIn_write_cmd_payload_address[31:0]               ), //i
    .io_push_payload_data        (io_gmbIn_write_cmd_payload_data[31:0]                  ), //i
    .io_push_payload_byteEnables (io_gmbIn_write_cmd_payload_byteEnables[3:0]            ), //i
    .io_push_payload_id          (io_gmbIn_write_cmd_payload_id[3:0]                     ), //i
    .io_push_payload_last        (io_gmbIn_write_cmd_payload_last                        ), //i
    .io_pop_valid                (io_gmbIn_write_cmd_fifo_io_pop_valid                   ), //o
    .io_pop_ready                (io_gmbIn_write_cmd_fifo_io_pop_fork_io_input_ready     ), //i
    .io_pop_payload_address      (io_gmbIn_write_cmd_fifo_io_pop_payload_address[31:0]   ), //o
    .io_pop_payload_data         (io_gmbIn_write_cmd_fifo_io_pop_payload_data[31:0]      ), //o
    .io_pop_payload_byteEnables  (io_gmbIn_write_cmd_fifo_io_pop_payload_byteEnables[3:0]), //o
    .io_pop_payload_id           (io_gmbIn_write_cmd_fifo_io_pop_payload_id[3:0]         ), //o
    .io_pop_payload_last         (io_gmbIn_write_cmd_fifo_io_pop_payload_last            ), //o
    .io_flush                    (1'b0                                                   ), //i
    .io_occupancy                (io_gmbIn_write_cmd_fifo_io_occupancy[1:0]              ), //o
    .io_availability             (io_gmbIn_write_cmd_fifo_io_availability[1:0]           ), //o
    .clk                         (clk                                                    ), //i
    .reset                       (reset                                                  )  //i
  );
  StreamFork io_gmbIn_write_cmd_fifo_io_pop_fork (
    .io_input_valid                   (io_gmbIn_write_cmd_fifo_io_pop_valid                                     ), //i
    .io_input_ready                   (io_gmbIn_write_cmd_fifo_io_pop_fork_io_input_ready                       ), //o
    .io_input_payload_address         (io_gmbIn_write_cmd_fifo_io_pop_payload_address[31:0]                     ), //i
    .io_input_payload_data            (io_gmbIn_write_cmd_fifo_io_pop_payload_data[31:0]                        ), //i
    .io_input_payload_byteEnables     (io_gmbIn_write_cmd_fifo_io_pop_payload_byteEnables[3:0]                  ), //i
    .io_input_payload_id              (io_gmbIn_write_cmd_fifo_io_pop_payload_id[3:0]                           ), //i
    .io_input_payload_last            (io_gmbIn_write_cmd_fifo_io_pop_payload_last                              ), //i
    .io_outputs_0_valid               (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_valid                   ), //o
    .io_outputs_0_ready               (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_ready        ), //i
    .io_outputs_0_payload_address     (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_address[31:0]   ), //o
    .io_outputs_0_payload_data        (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_data[31:0]      ), //o
    .io_outputs_0_payload_byteEnables (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_byteEnables[3:0]), //o
    .io_outputs_0_payload_id          (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_id[3:0]         ), //o
    .io_outputs_0_payload_last        (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_last            ), //o
    .io_outputs_1_valid               (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_valid                   ), //o
    .io_outputs_1_ready               (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_ready        ), //i
    .io_outputs_1_payload_address     (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_address[31:0]   ), //o
    .io_outputs_1_payload_data        (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_data[31:0]      ), //o
    .io_outputs_1_payload_byteEnables (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_byteEnables[3:0]), //o
    .io_outputs_1_payload_id          (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_id[3:0]         ), //o
    .io_outputs_1_payload_last        (io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_last            ), //o
    .clk                              (clk                                                                      ), //i
    .reset                            (reset                                                                    )  //i
  );
  StreamFifo_3 io_axiOut_b_fifo (
    .io_push_valid        (io_axiOut_b_valid                        ), //i
    .io_push_ready        (io_axiOut_b_fifo_io_push_ready           ), //o
    .io_push_payload_id   (io_axiOut_b_payload_id[3:0]              ), //i
    .io_push_payload_resp (io_axiOut_b_payload_resp[1:0]            ), //i
    .io_pop_valid         (io_axiOut_b_fifo_io_pop_valid            ), //o
    .io_pop_ready         (io_axiOut_b_fifo_io_pop_translated_ready ), //i
    .io_pop_payload_id    (io_axiOut_b_fifo_io_pop_payload_id[3:0]  ), //o
    .io_pop_payload_resp  (io_axiOut_b_fifo_io_pop_payload_resp[1:0]), //o
    .io_flush             (1'b0                                     ), //i
    .io_occupancy         (io_axiOut_b_fifo_io_occupancy[1:0]       ), //o
    .io_availability      (io_axiOut_b_fifo_io_availability[1:0]    ), //o
    .clk                  (clk                                      ), //i
    .reset                (reset                                    )  //i
  );
  assign io_gmbIn_read_cmd_ready = io_gmbIn_read_cmd_fifo_io_push_ready;
  assign io_gmbIn_read_cmd_fifo_io_pop_translated_valid = io_gmbIn_read_cmd_fifo_io_pop_valid;
  assign io_gmbIn_read_cmd_fifo_io_pop_translated_payload_addr = io_gmbIn_read_cmd_fifo_io_pop_payload_address;
  assign io_gmbIn_read_cmd_fifo_io_pop_translated_payload_id = io_gmbIn_read_cmd_fifo_io_pop_payload_id;
  assign io_gmbIn_read_cmd_fifo_io_pop_translated_payload_len = 8'h0;
  assign io_gmbIn_read_cmd_fifo_io_pop_translated_payload_size = 3'b010;
  assign io_gmbIn_read_cmd_fifo_io_pop_translated_payload_burst = 2'b01;
  assign io_axiOut_ar_valid = io_gmbIn_read_cmd_fifo_io_pop_translated_valid;
  assign io_gmbIn_read_cmd_fifo_io_pop_translated_ready = io_axiOut_ar_ready;
  assign io_axiOut_ar_payload_addr = io_gmbIn_read_cmd_fifo_io_pop_translated_payload_addr;
  assign io_axiOut_ar_payload_id = io_gmbIn_read_cmd_fifo_io_pop_translated_payload_id;
  assign io_axiOut_ar_payload_len = io_gmbIn_read_cmd_fifo_io_pop_translated_payload_len;
  assign io_axiOut_ar_payload_size = io_gmbIn_read_cmd_fifo_io_pop_translated_payload_size;
  assign io_axiOut_ar_payload_burst = io_gmbIn_read_cmd_fifo_io_pop_translated_payload_burst;
  assign io_axiOut_r_ready = io_axiOut_r_fifo_io_push_ready;
  assign io_axiOut_r_fifo_io_pop_translated_valid = io_axiOut_r_fifo_io_pop_valid;
  assign io_axiOut_r_fifo_io_pop_translated_payload_data = io_axiOut_r_fifo_io_pop_payload_data;
  assign io_axiOut_r_fifo_io_pop_translated_payload_error = (! (io_axiOut_r_fifo_io_pop_payload_resp == 2'b00));
  assign io_axiOut_r_fifo_io_pop_translated_payload_id = io_axiOut_r_fifo_io_pop_payload_id;
  assign io_gmbIn_read_rsp_valid = io_axiOut_r_fifo_io_pop_translated_valid;
  assign io_axiOut_r_fifo_io_pop_translated_ready = io_gmbIn_read_rsp_ready;
  assign io_gmbIn_read_rsp_payload_data = io_axiOut_r_fifo_io_pop_translated_payload_data;
  assign io_gmbIn_read_rsp_payload_error = io_axiOut_r_fifo_io_pop_translated_payload_error;
  assign io_gmbIn_read_rsp_payload_id = io_axiOut_r_fifo_io_pop_translated_payload_id;
  assign io_gmbIn_write_cmd_ready = io_gmbIn_write_cmd_fifo_io_push_ready;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_valid = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_valid;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_addr = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_address;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_id = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_payload_id;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_len = 8'h0;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_size = 3'b010;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_burst = 2'b01;
  assign io_axiOut_aw_valid = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_valid;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_ready = io_axiOut_aw_ready;
  assign io_axiOut_aw_payload_addr = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_addr;
  assign io_axiOut_aw_payload_id = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_id;
  assign io_axiOut_aw_payload_len = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_len;
  assign io_axiOut_aw_payload_size = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_size;
  assign io_axiOut_aw_payload_burst = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_0_translated_payload_burst;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_valid = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_valid;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_data = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_data;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_strb = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_payload_byteEnables;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_last = 1'b1;
  assign io_axiOut_w_valid = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_valid;
  assign io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_ready = io_axiOut_w_ready;
  assign io_axiOut_w_payload_data = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_data;
  assign io_axiOut_w_payload_strb = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_strb;
  assign io_axiOut_w_payload_last = io_gmbIn_write_cmd_fifo_io_pop_fork_io_outputs_1_translated_payload_last;
  assign io_axiOut_b_ready = io_axiOut_b_fifo_io_push_ready;
  assign io_axiOut_b_fifo_io_pop_translated_valid = io_axiOut_b_fifo_io_pop_valid;
  assign io_axiOut_b_fifo_io_pop_translated_payload_error = (! (io_axiOut_b_fifo_io_pop_payload_resp == 2'b00));
  assign io_axiOut_b_fifo_io_pop_translated_payload_id = io_axiOut_b_fifo_io_pop_payload_id;
  assign io_gmbIn_write_rsp_valid = io_axiOut_b_fifo_io_pop_translated_valid;
  assign io_axiOut_b_fifo_io_pop_translated_ready = io_gmbIn_write_rsp_ready;
  assign io_gmbIn_write_rsp_payload_error = io_axiOut_b_fifo_io_pop_translated_payload_error;
  assign io_gmbIn_write_rsp_payload_id = io_axiOut_b_fifo_io_pop_translated_payload_id;

endmodule

//InstructionPredecoder_3 replaced by InstructionPredecoder

//InstructionPredecoder_2 replaced by InstructionPredecoder

//InstructionPredecoder_1 replaced by InstructionPredecoder

module InstructionPredecoder (
  input  wire [31:0]   io_instruction,
  output reg           io_predecodeInfo_isBranch,
  output reg           io_predecodeInfo_isJump,
  output reg           io_predecodeInfo_isDirectJump,
  output reg  [31:0]   io_predecodeInfo_jumpOffset,
  output reg           io_predecodeInfo_isIdle,
  input  wire          clk,
  input  wire          reset
);

  wire       [27:0]   _zz_offset;
  wire       [5:0]    opcode;
  wire       [6:0]    opcode_7b;
  wire       [9:0]    idle_fixed_bits;
  wire       [25:0]   offs26;
  wire       [31:0]   offset;
  wire                when_InstructionPredecoder_l65;
  wire       [31:0]   _zz_1;

  assign _zz_offset = {offs26,2'b00};
  assign opcode = io_instruction[31 : 26];
  assign opcode_7b = io_instruction[31 : 25];
  assign idle_fixed_bits = io_instruction[24 : 15];
  always @(*) begin
    io_predecodeInfo_isBranch = 1'b0;
    case(opcode)
      6'h12, 6'h13, 6'h16, 6'h17, 6'h18, 6'h19, 6'h1a, 6'h1b : begin
        io_predecodeInfo_isBranch = 1'b1;
      end
      6'h14 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_predecodeInfo_isJump = 1'b0;
    case(opcode)
      6'h12, 6'h13, 6'h16, 6'h17, 6'h18, 6'h19, 6'h1a, 6'h1b : begin
      end
      6'h14 : begin
        io_predecodeInfo_isJump = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_predecodeInfo_isDirectJump = 1'b0;
    case(opcode)
      6'h12, 6'h13, 6'h16, 6'h17, 6'h18, 6'h19, 6'h1a, 6'h1b : begin
      end
      6'h14 : begin
        io_predecodeInfo_isDirectJump = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_predecodeInfo_jumpOffset = 32'h0;
    case(opcode)
      6'h12, 6'h13, 6'h16, 6'h17, 6'h18, 6'h19, 6'h1a, 6'h1b : begin
      end
      6'h14 : begin
        io_predecodeInfo_jumpOffset = offset;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_predecodeInfo_isIdle = 1'b0;
    if(when_InstructionPredecoder_l65) begin
      io_predecodeInfo_isIdle = 1'b1;
    end
  end

  assign offs26 = {io_instruction[25 : 16],io_instruction[15 : 0]};
  assign offset = {{4{_zz_offset[27]}}, _zz_offset};
  assign when_InstructionPredecoder_l65 = ((opcode_7b == 7'h03) && (idle_fixed_bits == 10'h091));
  assign _zz_1 = io_instruction;
  always @(posedge clk) begin
    if(reset) begin
    end else begin
      if(when_InstructionPredecoder_l65) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // InstructionPredecoder.scala:L67
          `else
            if(!1'b0) begin
              $display("NOTE(InstructionPredecoder.scala:67):  Found IDLE instruction: %x", _zz_1); // InstructionPredecoder.scala:L67
            end
          `endif
        `endif
      end
    end
  end


endmodule

module StreamFifo_12 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_pc,
  input  wire [31:0]   io_push_payload_instructions_0,
  input  wire [31:0]   io_push_payload_instructions_1,
  input  wire [31:0]   io_push_payload_instructions_2,
  input  wire [31:0]   io_push_payload_instructions_3,
  input  wire          io_push_payload_predecodeInfos_0_isBranch,
  input  wire          io_push_payload_predecodeInfos_0_isJump,
  input  wire          io_push_payload_predecodeInfos_0_isDirectJump,
  input  wire [31:0]   io_push_payload_predecodeInfos_0_jumpOffset,
  input  wire          io_push_payload_predecodeInfos_0_isIdle,
  input  wire          io_push_payload_predecodeInfos_1_isBranch,
  input  wire          io_push_payload_predecodeInfos_1_isJump,
  input  wire          io_push_payload_predecodeInfos_1_isDirectJump,
  input  wire [31:0]   io_push_payload_predecodeInfos_1_jumpOffset,
  input  wire          io_push_payload_predecodeInfos_1_isIdle,
  input  wire          io_push_payload_predecodeInfos_2_isBranch,
  input  wire          io_push_payload_predecodeInfos_2_isJump,
  input  wire          io_push_payload_predecodeInfos_2_isDirectJump,
  input  wire [31:0]   io_push_payload_predecodeInfos_2_jumpOffset,
  input  wire          io_push_payload_predecodeInfos_2_isIdle,
  input  wire          io_push_payload_predecodeInfos_3_isBranch,
  input  wire          io_push_payload_predecodeInfos_3_isJump,
  input  wire          io_push_payload_predecodeInfos_3_isDirectJump,
  input  wire [31:0]   io_push_payload_predecodeInfos_3_jumpOffset,
  input  wire          io_push_payload_predecodeInfos_3_isIdle,
  input  wire [3:0]    io_push_payload_branchMask,
  input  wire          io_push_payload_fault,
  input  wire [2:0]    io_push_payload_numValidInstructions,
  input  wire [1:0]    io_push_payload_startInstructionIndex,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_pc,
  output wire [31:0]   io_pop_payload_instructions_0,
  output wire [31:0]   io_pop_payload_instructions_1,
  output wire [31:0]   io_pop_payload_instructions_2,
  output wire [31:0]   io_pop_payload_instructions_3,
  output wire          io_pop_payload_predecodeInfos_0_isBranch,
  output wire          io_pop_payload_predecodeInfos_0_isJump,
  output wire          io_pop_payload_predecodeInfos_0_isDirectJump,
  output wire [31:0]   io_pop_payload_predecodeInfos_0_jumpOffset,
  output wire          io_pop_payload_predecodeInfos_0_isIdle,
  output wire          io_pop_payload_predecodeInfos_1_isBranch,
  output wire          io_pop_payload_predecodeInfos_1_isJump,
  output wire          io_pop_payload_predecodeInfos_1_isDirectJump,
  output wire [31:0]   io_pop_payload_predecodeInfos_1_jumpOffset,
  output wire          io_pop_payload_predecodeInfos_1_isIdle,
  output wire          io_pop_payload_predecodeInfos_2_isBranch,
  output wire          io_pop_payload_predecodeInfos_2_isJump,
  output wire          io_pop_payload_predecodeInfos_2_isDirectJump,
  output wire [31:0]   io_pop_payload_predecodeInfos_2_jumpOffset,
  output wire          io_pop_payload_predecodeInfos_2_isIdle,
  output wire          io_pop_payload_predecodeInfos_3_isBranch,
  output wire          io_pop_payload_predecodeInfos_3_isJump,
  output wire          io_pop_payload_predecodeInfos_3_isDirectJump,
  output wire [31:0]   io_pop_payload_predecodeInfos_3_jumpOffset,
  output wire          io_pop_payload_predecodeInfos_3_isIdle,
  output wire [3:0]    io_pop_payload_branchMask,
  output wire          io_pop_payload_fault,
  output wire [2:0]    io_pop_payload_numValidInstructions,
  output wire [1:0]    io_pop_payload_startInstructionIndex,
  input  wire          io_flush,
  output wire [1:0]    io_occupancy,
  output wire [1:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [313:0]  logic_ram_spinal_port1;
  wire       [313:0]  _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [1:0]    logic_ptr_push;
  reg        [1:0]    logic_ptr_pop;
  wire       [1:0]    logic_ptr_occupancy;
  wire       [1:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1455;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [0:0]    logic_push_onRam_write_payload_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_pc;
  wire       [31:0]   logic_push_onRam_write_payload_data_instructions_0;
  wire       [31:0]   logic_push_onRam_write_payload_data_instructions_1;
  wire       [31:0]   logic_push_onRam_write_payload_data_instructions_2;
  wire       [31:0]   logic_push_onRam_write_payload_data_instructions_3;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_0_isBranch;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_0_isJump;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_0_isDirectJump;
  wire       [31:0]   logic_push_onRam_write_payload_data_predecodeInfos_0_jumpOffset;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_0_isIdle;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_1_isBranch;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_1_isJump;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_1_isDirectJump;
  wire       [31:0]   logic_push_onRam_write_payload_data_predecodeInfos_1_jumpOffset;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_1_isIdle;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_2_isBranch;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_2_isJump;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_2_isDirectJump;
  wire       [31:0]   logic_push_onRam_write_payload_data_predecodeInfos_2_jumpOffset;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_2_isIdle;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_3_isBranch;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_3_isJump;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_3_isDirectJump;
  wire       [31:0]   logic_push_onRam_write_payload_data_predecodeInfos_3_jumpOffset;
  wire                logic_push_onRam_write_payload_data_predecodeInfos_3_isIdle;
  wire       [3:0]    logic_push_onRam_write_payload_data_branchMask;
  wire                logic_push_onRam_write_payload_data_fault;
  wire       [2:0]    logic_push_onRam_write_payload_data_numValidInstructions;
  wire       [1:0]    logic_push_onRam_write_payload_data_startInstructionIndex;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [0:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [0:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [0:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l477;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [0:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [31:0]   logic_pop_sync_readPort_rsp_pc;
  wire       [31:0]   logic_pop_sync_readPort_rsp_instructions_0;
  wire       [31:0]   logic_pop_sync_readPort_rsp_instructions_1;
  wire       [31:0]   logic_pop_sync_readPort_rsp_instructions_2;
  wire       [31:0]   logic_pop_sync_readPort_rsp_instructions_3;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_0_isJump;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_0_isDirectJump;
  wire       [31:0]   logic_pop_sync_readPort_rsp_predecodeInfos_0_jumpOffset;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_0_isIdle;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_1_isJump;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_1_isDirectJump;
  wire       [31:0]   logic_pop_sync_readPort_rsp_predecodeInfos_1_jumpOffset;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_1_isIdle;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_2_isJump;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_2_isDirectJump;
  wire       [31:0]   logic_pop_sync_readPort_rsp_predecodeInfos_2_jumpOffset;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_2_isIdle;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_3_isJump;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_3_isDirectJump;
  wire       [31:0]   logic_pop_sync_readPort_rsp_predecodeInfos_3_jumpOffset;
  wire                logic_pop_sync_readPort_rsp_predecodeInfos_3_isIdle;
  wire       [3:0]    logic_pop_sync_readPort_rsp_branchMask;
  wire                logic_pop_sync_readPort_rsp_fault;
  wire       [2:0]    logic_pop_sync_readPort_rsp_numValidInstructions;
  wire       [1:0]    logic_pop_sync_readPort_rsp_startInstructionIndex;
  wire       [313:0]  _zz_logic_pop_sync_readPort_rsp_pc;
  wire       [127:0]  _zz_logic_pop_sync_readPort_rsp_instructions_0;
  wire       [143:0]  _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch;
  wire       [35:0]   _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch_1;
  wire       [35:0]   _zz_logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch;
  wire       [35:0]   _zz_logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch;
  wire       [35:0]   _zz_logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch;
  wire                logic_pop_addressGen_toFlowFire_valid;
  wire       [0:0]    logic_pop_addressGen_toFlowFire_payload;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_pc;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_instructions_0;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_instructions_1;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_instructions_2;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_instructions_3;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isBranch;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isJump;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isDirectJump;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_jumpOffset;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isIdle;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isBranch;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isJump;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isDirectJump;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_jumpOffset;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isIdle;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isBranch;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isJump;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isDirectJump;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_jumpOffset;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isIdle;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isBranch;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isJump;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isDirectJump;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_jumpOffset;
  wire                logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isIdle;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_branchMask;
  wire                logic_pop_sync_readArbitation_translated_payload_fault;
  wire       [2:0]    logic_pop_sync_readArbitation_translated_payload_numValidInstructions;
  wire       [1:0]    logic_pop_sync_readArbitation_translated_payload_startInstructionIndex;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [1:0]    logic_pop_sync_popReg;
  (* ram_style = "block" *) reg [313:0] logic_ram [0:1];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_startInstructionIndex,{logic_push_onRam_write_payload_data_numValidInstructions,{logic_push_onRam_write_payload_data_fault,{logic_push_onRam_write_payload_data_branchMask,{{{logic_push_onRam_write_payload_data_predecodeInfos_3_isIdle,{logic_push_onRam_write_payload_data_predecodeInfos_3_jumpOffset,{logic_push_onRam_write_payload_data_predecodeInfos_3_isDirectJump,{logic_push_onRam_write_payload_data_predecodeInfos_3_isJump,logic_push_onRam_write_payload_data_predecodeInfos_3_isBranch}}}},{{logic_push_onRam_write_payload_data_predecodeInfos_2_isIdle,{logic_push_onRam_write_payload_data_predecodeInfos_2_jumpOffset,{logic_push_onRam_write_payload_data_predecodeInfos_2_isDirectJump,{logic_push_onRam_write_payload_data_predecodeInfos_2_isJump,logic_push_onRam_write_payload_data_predecodeInfos_2_isBranch}}}},{{logic_push_onRam_write_payload_data_predecodeInfos_1_isIdle,{logic_push_onRam_write_payload_data_predecodeInfos_1_jumpOffset,{logic_push_onRam_write_payload_data_predecodeInfos_1_isDirectJump,{logic_push_onRam_write_payload_data_predecodeInfos_1_isJump,logic_push_onRam_write_payload_data_predecodeInfos_1_isBranch}}}},{logic_push_onRam_write_payload_data_predecodeInfos_0_isIdle,{logic_push_onRam_write_payload_data_predecodeInfos_0_jumpOffset,{logic_push_onRam_write_payload_data_predecodeInfos_0_isDirectJump,{logic_push_onRam_write_payload_data_predecodeInfos_0_isJump,logic_push_onRam_write_payload_data_predecodeInfos_0_isBranch}}}}}}},{{logic_push_onRam_write_payload_data_instructions_3,{logic_push_onRam_write_payload_data_instructions_2,{logic_push_onRam_write_payload_data_instructions_1,logic_push_onRam_write_payload_data_instructions_0}}},logic_push_onRam_write_payload_data_pc}}}}}};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1455 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 2'b10) == 2'b00);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[0:0];
  assign logic_push_onRam_write_payload_data_pc = io_push_payload_pc;
  assign logic_push_onRam_write_payload_data_instructions_0 = io_push_payload_instructions_0;
  assign logic_push_onRam_write_payload_data_instructions_1 = io_push_payload_instructions_1;
  assign logic_push_onRam_write_payload_data_instructions_2 = io_push_payload_instructions_2;
  assign logic_push_onRam_write_payload_data_instructions_3 = io_push_payload_instructions_3;
  assign logic_push_onRam_write_payload_data_predecodeInfos_0_isBranch = io_push_payload_predecodeInfos_0_isBranch;
  assign logic_push_onRam_write_payload_data_predecodeInfos_0_isJump = io_push_payload_predecodeInfos_0_isJump;
  assign logic_push_onRam_write_payload_data_predecodeInfos_0_isDirectJump = io_push_payload_predecodeInfos_0_isDirectJump;
  assign logic_push_onRam_write_payload_data_predecodeInfos_0_jumpOffset = io_push_payload_predecodeInfos_0_jumpOffset;
  assign logic_push_onRam_write_payload_data_predecodeInfos_0_isIdle = io_push_payload_predecodeInfos_0_isIdle;
  assign logic_push_onRam_write_payload_data_predecodeInfos_1_isBranch = io_push_payload_predecodeInfos_1_isBranch;
  assign logic_push_onRam_write_payload_data_predecodeInfos_1_isJump = io_push_payload_predecodeInfos_1_isJump;
  assign logic_push_onRam_write_payload_data_predecodeInfos_1_isDirectJump = io_push_payload_predecodeInfos_1_isDirectJump;
  assign logic_push_onRam_write_payload_data_predecodeInfos_1_jumpOffset = io_push_payload_predecodeInfos_1_jumpOffset;
  assign logic_push_onRam_write_payload_data_predecodeInfos_1_isIdle = io_push_payload_predecodeInfos_1_isIdle;
  assign logic_push_onRam_write_payload_data_predecodeInfos_2_isBranch = io_push_payload_predecodeInfos_2_isBranch;
  assign logic_push_onRam_write_payload_data_predecodeInfos_2_isJump = io_push_payload_predecodeInfos_2_isJump;
  assign logic_push_onRam_write_payload_data_predecodeInfos_2_isDirectJump = io_push_payload_predecodeInfos_2_isDirectJump;
  assign logic_push_onRam_write_payload_data_predecodeInfos_2_jumpOffset = io_push_payload_predecodeInfos_2_jumpOffset;
  assign logic_push_onRam_write_payload_data_predecodeInfos_2_isIdle = io_push_payload_predecodeInfos_2_isIdle;
  assign logic_push_onRam_write_payload_data_predecodeInfos_3_isBranch = io_push_payload_predecodeInfos_3_isBranch;
  assign logic_push_onRam_write_payload_data_predecodeInfos_3_isJump = io_push_payload_predecodeInfos_3_isJump;
  assign logic_push_onRam_write_payload_data_predecodeInfos_3_isDirectJump = io_push_payload_predecodeInfos_3_isDirectJump;
  assign logic_push_onRam_write_payload_data_predecodeInfos_3_jumpOffset = io_push_payload_predecodeInfos_3_jumpOffset;
  assign logic_push_onRam_write_payload_data_predecodeInfos_3_isIdle = io_push_payload_predecodeInfos_3_isIdle;
  assign logic_push_onRam_write_payload_data_branchMask = io_push_payload_branchMask;
  assign logic_push_onRam_write_payload_data_fault = io_push_payload_fault;
  assign logic_push_onRam_write_payload_data_numValidInstructions = io_push_payload_numValidInstructions;
  assign logic_push_onRam_write_payload_data_startInstructionIndex = io_push_payload_startInstructionIndex;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[0:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l477) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_pc = logic_ram_spinal_port1;
  assign _zz_logic_pop_sync_readPort_rsp_instructions_0 = _zz_logic_pop_sync_readPort_rsp_pc[159 : 32];
  assign _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch = _zz_logic_pop_sync_readPort_rsp_pc[303 : 160];
  assign _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch_1 = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch[35 : 0];
  assign _zz_logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch[71 : 36];
  assign _zz_logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch[107 : 72];
  assign _zz_logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch[143 : 108];
  assign logic_pop_sync_readPort_rsp_pc = _zz_logic_pop_sync_readPort_rsp_pc[31 : 0];
  assign logic_pop_sync_readPort_rsp_instructions_0 = _zz_logic_pop_sync_readPort_rsp_instructions_0[31 : 0];
  assign logic_pop_sync_readPort_rsp_instructions_1 = _zz_logic_pop_sync_readPort_rsp_instructions_0[63 : 32];
  assign logic_pop_sync_readPort_rsp_instructions_2 = _zz_logic_pop_sync_readPort_rsp_instructions_0[95 : 64];
  assign logic_pop_sync_readPort_rsp_instructions_3 = _zz_logic_pop_sync_readPort_rsp_instructions_0[127 : 96];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch_1[0];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_0_isJump = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch_1[1];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_0_isDirectJump = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch_1[2];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_0_jumpOffset = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch_1[34 : 3];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_0_isIdle = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch_1[35];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch[0];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_1_isJump = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch[1];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_1_isDirectJump = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch[2];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_1_jumpOffset = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch[34 : 3];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_1_isIdle = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch[35];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch[0];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_2_isJump = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch[1];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_2_isDirectJump = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch[2];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_2_jumpOffset = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch[34 : 3];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_2_isIdle = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch[35];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch[0];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_3_isJump = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch[1];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_3_isDirectJump = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch[2];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_3_jumpOffset = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch[34 : 3];
  assign logic_pop_sync_readPort_rsp_predecodeInfos_3_isIdle = _zz_logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch[35];
  assign logic_pop_sync_readPort_rsp_branchMask = _zz_logic_pop_sync_readPort_rsp_pc[307 : 304];
  assign logic_pop_sync_readPort_rsp_fault = _zz_logic_pop_sync_readPort_rsp_pc[308];
  assign logic_pop_sync_readPort_rsp_numValidInstructions = _zz_logic_pop_sync_readPort_rsp_pc[311 : 309];
  assign logic_pop_sync_readPort_rsp_startInstructionIndex = _zz_logic_pop_sync_readPort_rsp_pc[313 : 312];
  assign logic_pop_addressGen_toFlowFire_valid = logic_pop_addressGen_fire;
  assign logic_pop_addressGen_toFlowFire_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_toFlowFire_valid;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_toFlowFire_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_pc = logic_pop_sync_readPort_rsp_pc;
  assign logic_pop_sync_readArbitation_translated_payload_instructions_0 = logic_pop_sync_readPort_rsp_instructions_0;
  assign logic_pop_sync_readArbitation_translated_payload_instructions_1 = logic_pop_sync_readPort_rsp_instructions_1;
  assign logic_pop_sync_readArbitation_translated_payload_instructions_2 = logic_pop_sync_readPort_rsp_instructions_2;
  assign logic_pop_sync_readArbitation_translated_payload_instructions_3 = logic_pop_sync_readPort_rsp_instructions_3;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isBranch = logic_pop_sync_readPort_rsp_predecodeInfos_0_isBranch;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isJump = logic_pop_sync_readPort_rsp_predecodeInfos_0_isJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isDirectJump = logic_pop_sync_readPort_rsp_predecodeInfos_0_isDirectJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_jumpOffset = logic_pop_sync_readPort_rsp_predecodeInfos_0_jumpOffset;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isIdle = logic_pop_sync_readPort_rsp_predecodeInfos_0_isIdle;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isBranch = logic_pop_sync_readPort_rsp_predecodeInfos_1_isBranch;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isJump = logic_pop_sync_readPort_rsp_predecodeInfos_1_isJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isDirectJump = logic_pop_sync_readPort_rsp_predecodeInfos_1_isDirectJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_jumpOffset = logic_pop_sync_readPort_rsp_predecodeInfos_1_jumpOffset;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isIdle = logic_pop_sync_readPort_rsp_predecodeInfos_1_isIdle;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isBranch = logic_pop_sync_readPort_rsp_predecodeInfos_2_isBranch;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isJump = logic_pop_sync_readPort_rsp_predecodeInfos_2_isJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isDirectJump = logic_pop_sync_readPort_rsp_predecodeInfos_2_isDirectJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_jumpOffset = logic_pop_sync_readPort_rsp_predecodeInfos_2_jumpOffset;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isIdle = logic_pop_sync_readPort_rsp_predecodeInfos_2_isIdle;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isBranch = logic_pop_sync_readPort_rsp_predecodeInfos_3_isBranch;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isJump = logic_pop_sync_readPort_rsp_predecodeInfos_3_isJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isDirectJump = logic_pop_sync_readPort_rsp_predecodeInfos_3_isDirectJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_jumpOffset = logic_pop_sync_readPort_rsp_predecodeInfos_3_jumpOffset;
  assign logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isIdle = logic_pop_sync_readPort_rsp_predecodeInfos_3_isIdle;
  assign logic_pop_sync_readArbitation_translated_payload_branchMask = logic_pop_sync_readPort_rsp_branchMask;
  assign logic_pop_sync_readArbitation_translated_payload_fault = logic_pop_sync_readPort_rsp_fault;
  assign logic_pop_sync_readArbitation_translated_payload_numValidInstructions = logic_pop_sync_readPort_rsp_numValidInstructions;
  assign logic_pop_sync_readArbitation_translated_payload_startInstructionIndex = logic_pop_sync_readPort_rsp_startInstructionIndex;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_pc = logic_pop_sync_readArbitation_translated_payload_pc;
  assign io_pop_payload_instructions_0 = logic_pop_sync_readArbitation_translated_payload_instructions_0;
  assign io_pop_payload_instructions_1 = logic_pop_sync_readArbitation_translated_payload_instructions_1;
  assign io_pop_payload_instructions_2 = logic_pop_sync_readArbitation_translated_payload_instructions_2;
  assign io_pop_payload_instructions_3 = logic_pop_sync_readArbitation_translated_payload_instructions_3;
  assign io_pop_payload_predecodeInfos_0_isBranch = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isBranch;
  assign io_pop_payload_predecodeInfos_0_isJump = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isJump;
  assign io_pop_payload_predecodeInfos_0_isDirectJump = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isDirectJump;
  assign io_pop_payload_predecodeInfos_0_jumpOffset = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_jumpOffset;
  assign io_pop_payload_predecodeInfos_0_isIdle = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_0_isIdle;
  assign io_pop_payload_predecodeInfos_1_isBranch = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isBranch;
  assign io_pop_payload_predecodeInfos_1_isJump = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isJump;
  assign io_pop_payload_predecodeInfos_1_isDirectJump = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isDirectJump;
  assign io_pop_payload_predecodeInfos_1_jumpOffset = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_jumpOffset;
  assign io_pop_payload_predecodeInfos_1_isIdle = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_1_isIdle;
  assign io_pop_payload_predecodeInfos_2_isBranch = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isBranch;
  assign io_pop_payload_predecodeInfos_2_isJump = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isJump;
  assign io_pop_payload_predecodeInfos_2_isDirectJump = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isDirectJump;
  assign io_pop_payload_predecodeInfos_2_jumpOffset = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_jumpOffset;
  assign io_pop_payload_predecodeInfos_2_isIdle = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_2_isIdle;
  assign io_pop_payload_predecodeInfos_3_isBranch = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isBranch;
  assign io_pop_payload_predecodeInfos_3_isJump = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isJump;
  assign io_pop_payload_predecodeInfos_3_isDirectJump = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isDirectJump;
  assign io_pop_payload_predecodeInfos_3_jumpOffset = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_jumpOffset;
  assign io_pop_payload_predecodeInfos_3_isIdle = logic_pop_sync_readArbitation_translated_payload_predecodeInfos_3_isIdle;
  assign io_pop_payload_branchMask = logic_pop_sync_readArbitation_translated_payload_branchMask;
  assign io_pop_payload_fault = logic_pop_sync_readArbitation_translated_payload_fault;
  assign io_pop_payload_numValidInstructions = logic_pop_sync_readArbitation_translated_payload_numValidInstructions;
  assign io_pop_payload_startInstructionIndex = logic_pop_sync_readArbitation_translated_payload_startInstructionIndex;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (2'b10 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 2'b00;
      logic_ptr_pop <= 2'b00;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 2'b00;
    end else begin
      if(when_Stream_l1455) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 2'b01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 2'b01);
      end
      if(io_flush) begin
        logic_ptr_push <= 2'b00;
        logic_ptr_pop <= 2'b00;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 2'b00;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module SmartDispatcher (
  input  wire          io_fetchGroupIn_valid,
  output wire          io_fetchGroupIn_ready,
  input  wire [31:0]   io_fetchGroupIn_payload_pc,
  input  wire [31:0]   io_fetchGroupIn_payload_instructions_0,
  input  wire [31:0]   io_fetchGroupIn_payload_instructions_1,
  input  wire [31:0]   io_fetchGroupIn_payload_instructions_2,
  input  wire [31:0]   io_fetchGroupIn_payload_instructions_3,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_0_isBranch,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_0_isJump,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_0_isDirectJump,
  input  wire [31:0]   io_fetchGroupIn_payload_predecodeInfos_0_jumpOffset,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_0_isIdle,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_1_isBranch,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_1_isJump,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_1_isDirectJump,
  input  wire [31:0]   io_fetchGroupIn_payload_predecodeInfos_1_jumpOffset,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_1_isIdle,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_2_isBranch,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_2_isJump,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_2_isDirectJump,
  input  wire [31:0]   io_fetchGroupIn_payload_predecodeInfos_2_jumpOffset,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_2_isIdle,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_3_isBranch,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_3_isJump,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_3_isDirectJump,
  input  wire [31:0]   io_fetchGroupIn_payload_predecodeInfos_3_jumpOffset,
  input  wire          io_fetchGroupIn_payload_predecodeInfos_3_isIdle,
  input  wire [3:0]    io_fetchGroupIn_payload_branchMask,
  input  wire          io_fetchGroupIn_payload_fault,
  input  wire [2:0]    io_fetchGroupIn_payload_numValidInstructions,
  input  wire [1:0]    io_fetchGroupIn_payload_startInstructionIndex,
  input  wire          io_bpuRsp_valid,
  input  wire          io_bpuRsp_payload_isTaken,
  input  wire [31:0]   io_bpuRsp_payload_target,
  input  wire [2:0]    io_bpuRsp_payload_transactionId,
  input  wire [31:0]   io_bpuRsp_payload_qPc,
  output reg           io_fetchOutput_valid,
  input  wire          io_fetchOutput_ready,
  output reg  [31:0]   io_fetchOutput_payload_pc,
  output reg  [31:0]   io_fetchOutput_payload_instruction,
  output reg           io_fetchOutput_payload_predecode_isBranch,
  output reg           io_fetchOutput_payload_predecode_isJump,
  output reg           io_fetchOutput_payload_predecode_isDirectJump,
  output reg  [31:0]   io_fetchOutput_payload_predecode_jumpOffset,
  output reg           io_fetchOutput_payload_predecode_isIdle,
  output reg           io_fetchOutput_payload_bpuPrediction_isTaken,
  output reg  [31:0]   io_fetchOutput_payload_bpuPrediction_target,
  output reg           io_fetchOutput_payload_bpuPrediction_wasPredicted,
  output reg           io_bpuQuery_valid,
  output reg  [31:0]   io_bpuQuery_payload_pc,
  output reg  [2:0]    io_bpuQuery_payload_transactionId,
  output reg           io_softRedirect_valid,
  output reg  [31:0]   io_softRedirect_payload,
  input  wire          io_flush,
  input  wire          clk,
  input  wire          reset
);
  localparam fsm_1_BOOT = 6'd1;
  localparam fsm_1_IDLE = 6'd2;
  localparam fsm_1_DISPATCHING = 6'd4;
  localparam fsm_1_WAITING_FOR_BPU = 6'd8;
  localparam fsm_1_SEND_BRANCH = 6'd16;
  localparam fsm_1_DRAINING_BPU = 6'd32;
  localparam fsm_1_BOOT_OH_ID = 0;
  localparam fsm_1_IDLE_OH_ID = 1;
  localparam fsm_1_DISPATCHING_OH_ID = 2;
  localparam fsm_1_WAITING_FOR_BPU_OH_ID = 3;
  localparam fsm_1_SEND_BRANCH_OH_ID = 4;
  localparam fsm_1_DRAINING_BPU_OH_ID = 5;

  wire       [31:0]   _zz_currentPcReg;
  reg        [31:0]   _zz_currentInstructionReg;
  reg                 _zz_currentPredecodeReg_isBranch;
  reg                 _zz_currentPredecodeReg_isJump;
  reg                 _zz_currentPredecodeReg_isDirectJump;
  reg        [31:0]   _zz_currentPredecodeReg_jumpOffset;
  reg                 _zz_currentPredecodeReg_isIdle;
  wire       [2:0]    _zz_lastInstructionIndexInGroup;
  wire       [2:0]    _zz_lastInstructionIndexInGroup_1;
  wire       [2:0]    _zz_isLastInstructionReg;
  reg                 _zz__zz_io_fetchOutput_payload_predecode_isBranch;
  reg                 _zz__zz_io_fetchOutput_payload_predecode_isJump;
  reg                 _zz__zz_io_fetchOutput_payload_predecode_isDirectJump;
  reg        [31:0]   _zz__zz_io_fetchOutput_payload_predecode_jumpOffset;
  reg                 _zz__zz_io_fetchOutput_payload_predecode_isIdle;
  wire       [31:0]   _zz__zz_io_fetchOutput_payload_pc;
  wire       [3:0]    _zz__zz_io_fetchOutput_payload_pc_1;
  reg        [31:0]   _zz__zz_io_fetchOutput_payload_instruction;
  wire       [2:0]    _zz_when_SmartDispatcher_l146;
  wire       [2:0]    _zz_when_SmartDispatcher_l146_1;
  wire       [31:0]   _zz_io_softRedirect_payload;
  reg        [31:0]   cycleReg;
  reg        [31:0]   fetchGroupReg_pc;
  reg        [31:0]   fetchGroupReg_instructions_0;
  reg        [31:0]   fetchGroupReg_instructions_1;
  reg        [31:0]   fetchGroupReg_instructions_2;
  reg        [31:0]   fetchGroupReg_instructions_3;
  reg                 fetchGroupReg_predecodeInfos_0_isBranch;
  reg                 fetchGroupReg_predecodeInfos_0_isJump;
  reg                 fetchGroupReg_predecodeInfos_0_isDirectJump;
  reg        [31:0]   fetchGroupReg_predecodeInfos_0_jumpOffset;
  reg                 fetchGroupReg_predecodeInfos_0_isIdle;
  reg                 fetchGroupReg_predecodeInfos_1_isBranch;
  reg                 fetchGroupReg_predecodeInfos_1_isJump;
  reg                 fetchGroupReg_predecodeInfos_1_isDirectJump;
  reg        [31:0]   fetchGroupReg_predecodeInfos_1_jumpOffset;
  reg                 fetchGroupReg_predecodeInfos_1_isIdle;
  reg                 fetchGroupReg_predecodeInfos_2_isBranch;
  reg                 fetchGroupReg_predecodeInfos_2_isJump;
  reg                 fetchGroupReg_predecodeInfos_2_isDirectJump;
  reg        [31:0]   fetchGroupReg_predecodeInfos_2_jumpOffset;
  reg                 fetchGroupReg_predecodeInfos_2_isIdle;
  reg                 fetchGroupReg_predecodeInfos_3_isBranch;
  reg                 fetchGroupReg_predecodeInfos_3_isJump;
  reg                 fetchGroupReg_predecodeInfos_3_isDirectJump;
  reg        [31:0]   fetchGroupReg_predecodeInfos_3_jumpOffset;
  reg                 fetchGroupReg_predecodeInfos_3_isIdle;
  reg        [3:0]    fetchGroupReg_branchMask;
  reg                 fetchGroupReg_fault;
  reg        [2:0]    fetchGroupReg_numValidInstructions;
  reg        [1:0]    fetchGroupReg_startInstructionIndex;
  reg                 isBusyReg;
  reg        [1:0]    dispatchIndexReg;
  reg        [2:0]    bpuInFlightCounterReg;
  reg        [2:0]    bpuTransIdCounterReg;
  reg        [31:0]   pendingBpuQueryReg_pc;
  reg        [31:0]   pendingBpuQueryReg_instruction;
  reg                 pendingBpuQueryReg_predecodeInfo_isBranch;
  reg                 pendingBpuQueryReg_predecodeInfo_isJump;
  reg                 pendingBpuQueryReg_predecodeInfo_isDirectJump;
  reg        [31:0]   pendingBpuQueryReg_predecodeInfo_jumpOffset;
  reg                 pendingBpuQueryReg_predecodeInfo_isIdle;
  reg        [2:0]    pendingBpuQueryReg_bpuTransactionId;
  reg        [31:0]   outputReg_pc;
  reg        [31:0]   outputReg_instruction;
  reg                 outputReg_predecode_isBranch;
  reg                 outputReg_predecode_isJump;
  reg                 outputReg_predecode_isDirectJump;
  reg        [31:0]   outputReg_predecode_jumpOffset;
  reg                 outputReg_predecode_isIdle;
  reg                 outputReg_bpuPrediction_isTaken;
  reg        [31:0]   outputReg_bpuPrediction_target;
  reg                 outputReg_bpuPrediction_wasPredicted;
  wire       [3:0]    pcIncrReg;
  wire       [31:0]   currentPcReg;
  wire       [31:0]   currentInstructionReg;
  wire                currentPredecodeReg_isBranch;
  wire                currentPredecodeReg_isJump;
  wire                currentPredecodeReg_isDirectJump;
  wire       [31:0]   currentPredecodeReg_jumpOffset;
  wire                currentPredecodeReg_isIdle;
  wire       [2:0]    lastInstructionIndexInGroup;
  wire                isLastInstructionReg;
  wire                hasValidInstructionReg;
  reg        [2:0]    fetchGroupReg_numValidInstructions_regNext;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg        [5:0]    fsm_stateReg;
  reg        [5:0]    fsm_stateNext;
  wire                when_SmartDispatcher_l108;
  wire                _zz_io_fetchOutput_payload_predecode_isBranch;
  wire                _zz_io_fetchOutput_payload_predecode_isJump;
  wire                _zz_io_fetchOutput_payload_predecode_isDirectJump;
  wire       [31:0]   _zz_io_fetchOutput_payload_predecode_jumpOffset;
  wire                _zz_io_fetchOutput_payload_predecode_isIdle;
  wire       [31:0]   _zz_io_fetchOutput_payload_pc;
  wire       [31:0]   _zz_io_fetchOutput_payload_instruction;
  wire                when_SmartDispatcher_l123;
  wire                when_SmartDispatcher_l146;
  wire                io_fetchGroupIn_fire;
  wire                when_SmartDispatcher_l206;
  wire                when_SmartDispatcher_l239;
  wire                when_SmartDispatcher_l279;
  wire                when_SmartDispatcher_l268;
  wire                when_SmartDispatcher_l273;
  wire                io_fetchOutput_fire;
  wire                when_SmartDispatcher_l316;
  wire                when_SmartDispatcher_l326;
  wire                when_SmartDispatcher_l347;
  wire                fsm_onExit_BOOT;
  wire                fsm_onExit_IDLE;
  wire                fsm_onExit_DISPATCHING;
  wire                fsm_onExit_WAITING_FOR_BPU;
  wire                fsm_onExit_SEND_BRANCH;
  wire                fsm_onExit_DRAINING_BPU;
  wire                fsm_onEntry_BOOT;
  wire                fsm_onEntry_IDLE;
  wire                fsm_onEntry_DISPATCHING;
  wire                fsm_onEntry_WAITING_FOR_BPU;
  wire                fsm_onEntry_SEND_BRANCH;
  wire                fsm_onEntry_DRAINING_BPU;
  reg        [2:0]    sim_fsmStateId;
  wire                when_SmartDispatcher_l381;
  wire                when_SmartDispatcher_l382;
  wire                when_SmartDispatcher_l383;
  wire                when_SmartDispatcher_l384;
  wire                when_SmartDispatcher_l385;
  `ifndef SYNTHESIS
  reg [119:0] fsm_stateReg_string;
  reg [119:0] fsm_stateNext_string;
  `endif


  assign _zz_currentPcReg = {28'd0, pcIncrReg};
  assign _zz_lastInstructionIndexInGroup = (_zz_lastInstructionIndexInGroup_1 + fetchGroupReg_numValidInstructions);
  assign _zz_lastInstructionIndexInGroup_1 = {1'd0, fetchGroupReg_startInstructionIndex};
  assign _zz_isLastInstructionReg = {1'd0, dispatchIndexReg};
  assign _zz__zz_io_fetchOutput_payload_pc_1 = ({2'd0,io_fetchGroupIn_payload_startInstructionIndex} <<< 2'd2);
  assign _zz__zz_io_fetchOutput_payload_pc = {28'd0, _zz__zz_io_fetchOutput_payload_pc_1};
  assign _zz_when_SmartDispatcher_l146 = {1'd0, io_fetchGroupIn_payload_startInstructionIndex};
  assign _zz_when_SmartDispatcher_l146_1 = (io_fetchGroupIn_payload_numValidInstructions - 3'b001);
  assign _zz_io_softRedirect_payload = (outputReg_pc + outputReg_predecode_jumpOffset);
  always @(*) begin
    case(dispatchIndexReg)
      2'b00 : begin
        _zz_currentInstructionReg = fetchGroupReg_instructions_0;
        _zz_currentPredecodeReg_isBranch = fetchGroupReg_predecodeInfos_0_isBranch;
        _zz_currentPredecodeReg_isJump = fetchGroupReg_predecodeInfos_0_isJump;
        _zz_currentPredecodeReg_isDirectJump = fetchGroupReg_predecodeInfos_0_isDirectJump;
        _zz_currentPredecodeReg_jumpOffset = fetchGroupReg_predecodeInfos_0_jumpOffset;
        _zz_currentPredecodeReg_isIdle = fetchGroupReg_predecodeInfos_0_isIdle;
      end
      2'b01 : begin
        _zz_currentInstructionReg = fetchGroupReg_instructions_1;
        _zz_currentPredecodeReg_isBranch = fetchGroupReg_predecodeInfos_1_isBranch;
        _zz_currentPredecodeReg_isJump = fetchGroupReg_predecodeInfos_1_isJump;
        _zz_currentPredecodeReg_isDirectJump = fetchGroupReg_predecodeInfos_1_isDirectJump;
        _zz_currentPredecodeReg_jumpOffset = fetchGroupReg_predecodeInfos_1_jumpOffset;
        _zz_currentPredecodeReg_isIdle = fetchGroupReg_predecodeInfos_1_isIdle;
      end
      2'b10 : begin
        _zz_currentInstructionReg = fetchGroupReg_instructions_2;
        _zz_currentPredecodeReg_isBranch = fetchGroupReg_predecodeInfos_2_isBranch;
        _zz_currentPredecodeReg_isJump = fetchGroupReg_predecodeInfos_2_isJump;
        _zz_currentPredecodeReg_isDirectJump = fetchGroupReg_predecodeInfos_2_isDirectJump;
        _zz_currentPredecodeReg_jumpOffset = fetchGroupReg_predecodeInfos_2_jumpOffset;
        _zz_currentPredecodeReg_isIdle = fetchGroupReg_predecodeInfos_2_isIdle;
      end
      default : begin
        _zz_currentInstructionReg = fetchGroupReg_instructions_3;
        _zz_currentPredecodeReg_isBranch = fetchGroupReg_predecodeInfos_3_isBranch;
        _zz_currentPredecodeReg_isJump = fetchGroupReg_predecodeInfos_3_isJump;
        _zz_currentPredecodeReg_isDirectJump = fetchGroupReg_predecodeInfos_3_isDirectJump;
        _zz_currentPredecodeReg_jumpOffset = fetchGroupReg_predecodeInfos_3_jumpOffset;
        _zz_currentPredecodeReg_isIdle = fetchGroupReg_predecodeInfos_3_isIdle;
      end
    endcase
  end

  always @(*) begin
    case(io_fetchGroupIn_payload_startInstructionIndex)
      2'b00 : begin
        _zz__zz_io_fetchOutput_payload_predecode_isBranch = io_fetchGroupIn_payload_predecodeInfos_0_isBranch;
        _zz__zz_io_fetchOutput_payload_predecode_isJump = io_fetchGroupIn_payload_predecodeInfos_0_isJump;
        _zz__zz_io_fetchOutput_payload_predecode_isDirectJump = io_fetchGroupIn_payload_predecodeInfos_0_isDirectJump;
        _zz__zz_io_fetchOutput_payload_predecode_jumpOffset = io_fetchGroupIn_payload_predecodeInfos_0_jumpOffset;
        _zz__zz_io_fetchOutput_payload_predecode_isIdle = io_fetchGroupIn_payload_predecodeInfos_0_isIdle;
        _zz__zz_io_fetchOutput_payload_instruction = io_fetchGroupIn_payload_instructions_0;
      end
      2'b01 : begin
        _zz__zz_io_fetchOutput_payload_predecode_isBranch = io_fetchGroupIn_payload_predecodeInfos_1_isBranch;
        _zz__zz_io_fetchOutput_payload_predecode_isJump = io_fetchGroupIn_payload_predecodeInfos_1_isJump;
        _zz__zz_io_fetchOutput_payload_predecode_isDirectJump = io_fetchGroupIn_payload_predecodeInfos_1_isDirectJump;
        _zz__zz_io_fetchOutput_payload_predecode_jumpOffset = io_fetchGroupIn_payload_predecodeInfos_1_jumpOffset;
        _zz__zz_io_fetchOutput_payload_predecode_isIdle = io_fetchGroupIn_payload_predecodeInfos_1_isIdle;
        _zz__zz_io_fetchOutput_payload_instruction = io_fetchGroupIn_payload_instructions_1;
      end
      2'b10 : begin
        _zz__zz_io_fetchOutput_payload_predecode_isBranch = io_fetchGroupIn_payload_predecodeInfos_2_isBranch;
        _zz__zz_io_fetchOutput_payload_predecode_isJump = io_fetchGroupIn_payload_predecodeInfos_2_isJump;
        _zz__zz_io_fetchOutput_payload_predecode_isDirectJump = io_fetchGroupIn_payload_predecodeInfos_2_isDirectJump;
        _zz__zz_io_fetchOutput_payload_predecode_jumpOffset = io_fetchGroupIn_payload_predecodeInfos_2_jumpOffset;
        _zz__zz_io_fetchOutput_payload_predecode_isIdle = io_fetchGroupIn_payload_predecodeInfos_2_isIdle;
        _zz__zz_io_fetchOutput_payload_instruction = io_fetchGroupIn_payload_instructions_2;
      end
      default : begin
        _zz__zz_io_fetchOutput_payload_predecode_isBranch = io_fetchGroupIn_payload_predecodeInfos_3_isBranch;
        _zz__zz_io_fetchOutput_payload_predecode_isJump = io_fetchGroupIn_payload_predecodeInfos_3_isJump;
        _zz__zz_io_fetchOutput_payload_predecode_isDirectJump = io_fetchGroupIn_payload_predecodeInfos_3_isDirectJump;
        _zz__zz_io_fetchOutput_payload_predecode_jumpOffset = io_fetchGroupIn_payload_predecodeInfos_3_jumpOffset;
        _zz__zz_io_fetchOutput_payload_predecode_isIdle = io_fetchGroupIn_payload_predecodeInfos_3_isIdle;
        _zz__zz_io_fetchOutput_payload_instruction = io_fetchGroupIn_payload_instructions_3;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_1_BOOT : fsm_stateReg_string = "BOOT           ";
      fsm_1_IDLE : fsm_stateReg_string = "IDLE           ";
      fsm_1_DISPATCHING : fsm_stateReg_string = "DISPATCHING    ";
      fsm_1_WAITING_FOR_BPU : fsm_stateReg_string = "WAITING_FOR_BPU";
      fsm_1_SEND_BRANCH : fsm_stateReg_string = "SEND_BRANCH    ";
      fsm_1_DRAINING_BPU : fsm_stateReg_string = "DRAINING_BPU   ";
      default : fsm_stateReg_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_1_BOOT : fsm_stateNext_string = "BOOT           ";
      fsm_1_IDLE : fsm_stateNext_string = "IDLE           ";
      fsm_1_DISPATCHING : fsm_stateNext_string = "DISPATCHING    ";
      fsm_1_WAITING_FOR_BPU : fsm_stateNext_string = "WAITING_FOR_BPU";
      fsm_1_SEND_BRANCH : fsm_stateNext_string = "SEND_BRANCH    ";
      fsm_1_DRAINING_BPU : fsm_stateNext_string = "DRAINING_BPU   ";
      default : fsm_stateNext_string = "???????????????";
    endcase
  end
  `endif

  always @(*) begin
    io_fetchOutput_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_valid = 1'b1;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_valid = 1'b1;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_valid = 1'b1;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_pc = _zz_io_fetchOutput_payload_pc;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_pc = currentPcReg;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_pc = outputReg_pc;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_instruction = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_instruction = _zz_io_fetchOutput_payload_instruction;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_instruction = currentInstructionReg;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_instruction = outputReg_instruction;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_predecode_isBranch = 1'bx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_predecode_isBranch = _zz_io_fetchOutput_payload_predecode_isBranch;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_predecode_isBranch = currentPredecodeReg_isBranch;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_predecode_isBranch = outputReg_predecode_isBranch;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_predecode_isJump = 1'bx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_predecode_isJump = _zz_io_fetchOutput_payload_predecode_isJump;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_predecode_isJump = currentPredecodeReg_isJump;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_predecode_isJump = outputReg_predecode_isJump;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_predecode_isDirectJump = 1'bx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_predecode_isDirectJump = _zz_io_fetchOutput_payload_predecode_isDirectJump;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_predecode_isDirectJump = currentPredecodeReg_isDirectJump;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_predecode_isDirectJump = outputReg_predecode_isDirectJump;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_predecode_jumpOffset = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_predecode_jumpOffset = _zz_io_fetchOutput_payload_predecode_jumpOffset;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_predecode_jumpOffset = currentPredecodeReg_jumpOffset;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_predecode_jumpOffset = outputReg_predecode_jumpOffset;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_predecode_isIdle = 1'bx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_predecode_isIdle = _zz_io_fetchOutput_payload_predecode_isIdle;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_predecode_isIdle = currentPredecodeReg_isIdle;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_predecode_isIdle = outputReg_predecode_isIdle;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_bpuPrediction_isTaken = 1'bx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_bpuPrediction_isTaken = 1'b0;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_bpuPrediction_isTaken = 1'b0;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_bpuPrediction_isTaken = outputReg_bpuPrediction_isTaken;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_bpuPrediction_target = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_bpuPrediction_target = 32'h0;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_bpuPrediction_target = 32'h0;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_bpuPrediction_target = outputReg_bpuPrediction_target;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_fetchOutput_payload_bpuPrediction_wasPredicted = 1'bx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                io_fetchOutput_payload_bpuPrediction_wasPredicted = 1'b0;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                io_fetchOutput_payload_bpuPrediction_wasPredicted = 1'b0;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          io_fetchOutput_payload_bpuPrediction_wasPredicted = outputReg_bpuPrediction_wasPredicted;
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_bpuQuery_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(!when_SmartDispatcher_l123) begin
                io_bpuQuery_valid = 1'b1;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(when_SmartDispatcher_l206) begin
                io_bpuQuery_valid = 1'b1;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_bpuQuery_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(!when_SmartDispatcher_l123) begin
                io_bpuQuery_payload_pc = _zz_io_fetchOutput_payload_pc;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(when_SmartDispatcher_l206) begin
                io_bpuQuery_payload_pc = currentPcReg;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_bpuQuery_payload_transactionId = 3'bxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(!when_SmartDispatcher_l123) begin
                io_bpuQuery_payload_transactionId = bpuTransIdCounterReg;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(when_SmartDispatcher_l206) begin
                io_bpuQuery_payload_transactionId = bpuTransIdCounterReg;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_softRedirect_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                if(io_fetchOutput_ready) begin
                  if(_zz_io_fetchOutput_payload_predecode_isDirectJump) begin
                    io_softRedirect_valid = 1'b1;
                  end
                end
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                if(io_fetchOutput_ready) begin
                  if(currentPredecodeReg_isDirectJump) begin
                    io_softRedirect_valid = 1'b1;
                  end
                end
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchOutput_fire) begin
            if(when_SmartDispatcher_l316) begin
              io_softRedirect_valid = 1'b1;
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_softRedirect_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                if(io_fetchOutput_ready) begin
                  if(_zz_io_fetchOutput_payload_predecode_isDirectJump) begin
                    io_softRedirect_payload = (_zz_io_fetchOutput_payload_pc + _zz_io_fetchOutput_payload_predecode_jumpOffset);
                  end
                end
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(!when_SmartDispatcher_l206) begin
                if(io_fetchOutput_ready) begin
                  if(currentPredecodeReg_isDirectJump) begin
                    io_softRedirect_payload = (currentPcReg + currentPredecodeReg_jumpOffset);
                  end
                end
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchOutput_fire) begin
            if(when_SmartDispatcher_l316) begin
              io_softRedirect_payload = (outputReg_predecode_isDirectJump ? _zz_io_softRedirect_payload : outputReg_bpuPrediction_target);
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign io_fetchGroupIn_ready = (! isBusyReg);
  assign pcIncrReg = ({2'd0,dispatchIndexReg} <<< 2'd2);
  assign currentPcReg = (fetchGroupReg_pc + _zz_currentPcReg);
  assign currentInstructionReg = _zz_currentInstructionReg;
  assign currentPredecodeReg_isBranch = _zz_currentPredecodeReg_isBranch;
  assign currentPredecodeReg_isJump = _zz_currentPredecodeReg_isJump;
  assign currentPredecodeReg_isDirectJump = _zz_currentPredecodeReg_isDirectJump;
  assign currentPredecodeReg_jumpOffset = _zz_currentPredecodeReg_jumpOffset;
  assign currentPredecodeReg_isIdle = _zz_currentPredecodeReg_isIdle;
  assign lastInstructionIndexInGroup = (_zz_lastInstructionIndexInGroup - 3'b001);
  assign isLastInstructionReg = (_zz_isLastInstructionReg == lastInstructionIndexInGroup);
  assign hasValidInstructionReg = (3'b000 < fetchGroupReg_numValidInstructions);
  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(io_flush) begin
          fsm_stateNext = fsm_1_IDLE;
        end else begin
          if(io_fetchGroupIn_fire) begin
            if(when_SmartDispatcher_l108) begin
              fsm_stateNext = fsm_1_IDLE;
            end else begin
              if(when_SmartDispatcher_l123) begin
                if(io_fetchOutput_ready) begin
                  if(_zz_io_fetchOutput_payload_predecode_isDirectJump) begin
                    fsm_stateNext = fsm_1_IDLE;
                  end else begin
                    if(when_SmartDispatcher_l146) begin
                      fsm_stateNext = fsm_1_IDLE;
                    end else begin
                      fsm_stateNext = fsm_1_DISPATCHING;
                    end
                  end
                end else begin
                  fsm_stateNext = fsm_1_SEND_BRANCH;
                end
              end else begin
                fsm_stateNext = fsm_1_WAITING_FOR_BPU;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(io_flush) begin
          fsm_stateNext = fsm_1_DRAINING_BPU;
        end else begin
          if(isBusyReg) begin
            if(fetchGroupReg_fault) begin
              fsm_stateNext = fsm_1_IDLE;
            end else begin
              if(when_SmartDispatcher_l206) begin
                fsm_stateNext = fsm_1_WAITING_FOR_BPU;
              end else begin
                if(io_fetchOutput_ready) begin
                  if(when_SmartDispatcher_l239) begin
                    fsm_stateNext = fsm_1_IDLE;
                  end
                end
              end
            end
          end else begin
            fsm_stateNext = fsm_1_IDLE;
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
        if(io_flush) begin
          fsm_stateNext = fsm_1_DRAINING_BPU;
        end else begin
          if(when_SmartDispatcher_l279) begin
            fsm_stateNext = fsm_1_SEND_BRANCH;
          end
        end
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
        if(io_flush) begin
          fsm_stateNext = fsm_1_DRAINING_BPU;
        end else begin
          if(io_fetchOutput_fire) begin
            if(when_SmartDispatcher_l326) begin
              fsm_stateNext = fsm_1_IDLE;
            end else begin
              fsm_stateNext = fsm_1_DISPATCHING;
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
        if(when_SmartDispatcher_l347) begin
          fsm_stateNext = fsm_1_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_1_IDLE;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_1_BOOT;
    end
  end

  assign when_SmartDispatcher_l108 = (io_fetchGroupIn_payload_numValidInstructions == 3'b000);
  assign _zz_io_fetchOutput_payload_predecode_isBranch = _zz__zz_io_fetchOutput_payload_predecode_isBranch;
  assign _zz_io_fetchOutput_payload_predecode_isJump = _zz__zz_io_fetchOutput_payload_predecode_isJump;
  assign _zz_io_fetchOutput_payload_predecode_isDirectJump = _zz__zz_io_fetchOutput_payload_predecode_isDirectJump;
  assign _zz_io_fetchOutput_payload_predecode_jumpOffset = _zz__zz_io_fetchOutput_payload_predecode_jumpOffset;
  assign _zz_io_fetchOutput_payload_predecode_isIdle = _zz__zz_io_fetchOutput_payload_predecode_isIdle;
  assign _zz_io_fetchOutput_payload_pc = (io_fetchGroupIn_payload_pc + _zz__zz_io_fetchOutput_payload_pc);
  assign _zz_io_fetchOutput_payload_instruction = _zz__zz_io_fetchOutput_payload_instruction;
  assign when_SmartDispatcher_l123 = (! _zz_io_fetchOutput_payload_predecode_isBranch);
  assign when_SmartDispatcher_l146 = (_zz_when_SmartDispatcher_l146 == _zz_when_SmartDispatcher_l146_1);
  assign io_fetchGroupIn_fire = (io_fetchGroupIn_valid && io_fetchGroupIn_ready);
  assign when_SmartDispatcher_l206 = (currentPredecodeReg_isBranch && (! currentPredecodeReg_isDirectJump));
  assign when_SmartDispatcher_l239 = (isLastInstructionReg || currentPredecodeReg_isDirectJump);
  assign when_SmartDispatcher_l279 = (io_bpuRsp_valid && (io_bpuRsp_payload_transactionId == pendingBpuQueryReg_bpuTransactionId));
  assign when_SmartDispatcher_l268 = (! when_SmartDispatcher_l279);
  assign when_SmartDispatcher_l273 = (isBusyReg && (! when_SmartDispatcher_l279));
  assign io_fetchOutput_fire = (io_fetchOutput_valid && io_fetchOutput_ready);
  assign when_SmartDispatcher_l316 = (outputReg_predecode_isDirectJump || (outputReg_bpuPrediction_wasPredicted && outputReg_bpuPrediction_isTaken));
  assign when_SmartDispatcher_l326 = (isLastInstructionReg || when_SmartDispatcher_l316);
  assign when_SmartDispatcher_l347 = (bpuInFlightCounterReg == 3'b000);
  assign fsm_onExit_BOOT = ((! fsm_stateNext[fsm_1_BOOT_OH_ID]) && (fsm_stateReg[fsm_1_BOOT_OH_ID]));
  assign fsm_onExit_IDLE = ((! fsm_stateNext[fsm_1_IDLE_OH_ID]) && (fsm_stateReg[fsm_1_IDLE_OH_ID]));
  assign fsm_onExit_DISPATCHING = ((! fsm_stateNext[fsm_1_DISPATCHING_OH_ID]) && (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]));
  assign fsm_onExit_WAITING_FOR_BPU = ((! fsm_stateNext[fsm_1_WAITING_FOR_BPU_OH_ID]) && (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]));
  assign fsm_onExit_SEND_BRANCH = ((! fsm_stateNext[fsm_1_SEND_BRANCH_OH_ID]) && (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]));
  assign fsm_onExit_DRAINING_BPU = ((! fsm_stateNext[fsm_1_DRAINING_BPU_OH_ID]) && (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]));
  assign fsm_onEntry_BOOT = ((fsm_stateNext[fsm_1_BOOT_OH_ID]) && (! fsm_stateReg[fsm_1_BOOT_OH_ID]));
  assign fsm_onEntry_IDLE = ((fsm_stateNext[fsm_1_IDLE_OH_ID]) && (! fsm_stateReg[fsm_1_IDLE_OH_ID]));
  assign fsm_onEntry_DISPATCHING = ((fsm_stateNext[fsm_1_DISPATCHING_OH_ID]) && (! fsm_stateReg[fsm_1_DISPATCHING_OH_ID]));
  assign fsm_onEntry_WAITING_FOR_BPU = ((fsm_stateNext[fsm_1_WAITING_FOR_BPU_OH_ID]) && (! fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]));
  assign fsm_onEntry_SEND_BRANCH = ((fsm_stateNext[fsm_1_SEND_BRANCH_OH_ID]) && (! fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]));
  assign fsm_onEntry_DRAINING_BPU = ((fsm_stateNext[fsm_1_DRAINING_BPU_OH_ID]) && (! fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]));
  assign when_SmartDispatcher_l381 = (fsm_stateReg[fsm_1_IDLE_OH_ID]);
  always @(*) begin
    if(when_SmartDispatcher_l381) begin
      sim_fsmStateId = 3'b000;
    end else begin
      if(when_SmartDispatcher_l382) begin
        sim_fsmStateId = 3'b001;
      end else begin
        if(when_SmartDispatcher_l383) begin
          sim_fsmStateId = 3'b010;
        end else begin
          if(when_SmartDispatcher_l384) begin
            sim_fsmStateId = 3'b011;
          end else begin
            if(when_SmartDispatcher_l385) begin
              sim_fsmStateId = 3'b100;
            end else begin
              sim_fsmStateId = 3'b101;
            end
          end
        end
      end
    end
  end

  assign when_SmartDispatcher_l382 = (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]);
  assign when_SmartDispatcher_l383 = (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]);
  assign when_SmartDispatcher_l384 = (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]);
  assign when_SmartDispatcher_l385 = (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]);
  always @(posedge clk) begin
    if(reset) begin
      cycleReg <= 32'h0;
      isBusyReg <= 1'b0;
      dispatchIndexReg <= 2'b00;
      bpuInFlightCounterReg <= 3'b000;
      bpuTransIdCounterReg <= 3'b000;
      fetchGroupReg_numValidInstructions_regNext <= 3'b000;
      fsm_stateReg <= fsm_1_BOOT;
    end else begin
      cycleReg <= (cycleReg + 32'h00000001);
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // SmartDispatcher.scala:L25
        `else
          if(!1'b0) begin
            $display("NOTE(SmartDispatcher.scala:25):  ------ RAW INSTR DISPATCHER CYCLE: %x", cycleReg); // SmartDispatcher.scala:L25
          end
        `endif
      `endif
      fetchGroupReg_numValidInstructions_regNext <= fetchGroupReg_numValidInstructions;
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // SmartDispatcher.scala:L57
        `else
          if(!1'b0) begin
            $display("NOTE(SmartDispatcher.scala:57):    DEBUG-VALID: fetchGroupReg numValidInstructions is %x, last cycle it is %x", fetchGroupReg_numValidInstructions, fetchGroupReg_numValidInstructions_regNext); // SmartDispatcher.scala:L57
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // SmartDispatcher.scala:L58
        `else
          if(!1'b0) begin
            $display("NOTE(SmartDispatcher.scala:58):    DEBUG: currentPc=0x%x, currentInstructionReg=0x%x, currentPredecodeReg.isBranch=%x, currentPredecodeReg.isDirectJump=%x", currentPcReg, currentInstructionReg, currentPredecodeReg_isBranch, currentPredecodeReg_isDirectJump); // SmartDispatcher.scala:L58
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // SmartDispatcher.scala:L59
        `else
          if(!1'b0) begin
            $display("NOTE(SmartDispatcher.scala:59):    DEBUG: fetchGroupReg.numValidInstructions=%x, dispatchIndexReg=%x", fetchGroupReg_numValidInstructions, dispatchIndexReg); // SmartDispatcher.scala:L59
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // SmartDispatcher.scala:L60
        `else
          if(!1'b0) begin
            $display("NOTE(SmartDispatcher.scala:60):    DEBUG: isLastInstruction=%x", isLastInstructionReg); // SmartDispatcher.scala:L60
          end
        `endif
      `endif
      if(io_bpuQuery_valid) begin
        bpuInFlightCounterReg <= (bpuInFlightCounterReg + 3'b001);
        bpuTransIdCounterReg <= (bpuTransIdCounterReg + 3'b001);
      end
      if(io_bpuRsp_valid) begin
        bpuInFlightCounterReg <= (bpuInFlightCounterReg - 3'b001);
      end
      fsm_stateReg <= fsm_stateNext;
      (* parallel_case *)
      case(1) // synthesis parallel_case
        (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
          if(io_flush) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // SmartDispatcher.scala:L88
              `else
                if(!1'b0) begin
                  $display("NOTE(SmartDispatcher.scala:88):  DISPATCHER-IDLE: Flush asserted, remaining in IDLE."); // SmartDispatcher.scala:L88
                end
              `endif
            `endif
          end else begin
            if(io_fetchGroupIn_fire) begin
              isBusyReg <= 1'b1;
              dispatchIndexReg <= io_fetchGroupIn_payload_startInstructionIndex;
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L99
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:99):    DEBUG-ASSIGN: dispatchIndexReg assigned 0 from IDLE"); // SmartDispatcher.scala:L99
                  end
                `endif
              `endif
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L103
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:103):  DISPATCHER-IDLE: New Group Received. PC=0x%x.", io_fetchGroupIn_payload_pc); // SmartDispatcher.scala:L103
                  end
                `endif
              `endif
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L104
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:104):    DEBUG-IDLE-LOAD-PAYLOAD: io.fetchGroupIn.payload.numValidInstructions=%x", io_fetchGroupIn_payload_numValidInstructions); // SmartDispatcher.scala:L104
                  end
                `endif
              `endif
              if(when_SmartDispatcher_l108) begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // SmartDispatcher.scala:L109
                  `else
                    if(!1'b0) begin
                      $display("NOTE(SmartDispatcher.scala:109):  DISPATCHER-IDLE: Received empty FetchGroup (numValidInstructions=0). Going back to IDLE."); // SmartDispatcher.scala:L109
                    end
                  `endif
                `endif
                isBusyReg <= 1'b0;
                dispatchIndexReg <= 2'b00;
              end else begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // SmartDispatcher.scala:L120
                  `else
                    if(!1'b0) begin
                      $display("NOTE(SmartDispatcher.scala:120):  DISPATCHER-IDLE: Analyzing first instruction (PC=0x%x, isBranch=%x).", _zz_io_fetchOutput_payload_pc, _zz_io_fetchOutput_payload_predecode_isBranch); // SmartDispatcher.scala:L120
                    end
                  `endif
                `endif
                if(when_SmartDispatcher_l123) begin
                  `ifndef SYNTHESIS
                    `ifdef FORMAL
                      assert(1'b0); // SmartDispatcher.scala:L124
                    `else
                      if(!1'b0) begin
                        $display("NOTE(SmartDispatcher.scala:124):  DISPATCHER-IDLE: First instruction is Fast Path. PC=0x%x", _zz_io_fetchOutput_payload_pc); // SmartDispatcher.scala:L124
                      end
                    `endif
                  `endif
                  if(io_fetchOutput_ready) begin
                    `ifndef SYNTHESIS
                      `ifdef FORMAL
                        assert(1'b0); // SmartDispatcher.scala:L133
                      `else
                        if(!1'b0) begin
                          $display("NOTE(SmartDispatcher.scala:133):  DISPATCHER-IDLE: First instruction (fast path) fired."); // SmartDispatcher.scala:L133
                        end
                      `endif
                    `endif
                    if(_zz_io_fetchOutput_payload_predecode_isDirectJump) begin
                      `ifndef SYNTHESIS
                        `ifdef FORMAL
                          assert(1'b0); // SmartDispatcher.scala:L137
                        `else
                          if(!1'b0) begin
                            $display("NOTE(SmartDispatcher.scala:137):  DISPATCHER-IDLE: First instruction is a direct jump. Redirecting to 0x%x.", io_softRedirect_payload); // SmartDispatcher.scala:L137
                          end
                        `endif
                      `endif
                      dispatchIndexReg <= 2'b00;
                      isBusyReg <= 1'b0;
                    end else begin
                      `ifndef SYNTHESIS
                        `ifdef FORMAL
                          assert(1'b0); // SmartDispatcher.scala:L144
                        `else
                          if(!1'b0) begin
                            $display("NOTE(SmartDispatcher.scala:144):    DEBUG-IDLE-FIRST-ISLAST: fetchGroupReg.numValidInstructions=%x, isFirstInstructionLast=%x", fetchGroupReg_numValidInstructions, when_SmartDispatcher_l146); // SmartDispatcher.scala:L144
                          end
                        `endif
                      `endif
                      if(when_SmartDispatcher_l146) begin
                        `ifndef SYNTHESIS
                          `ifdef FORMAL
                            assert(1'b0); // SmartDispatcher.scala:L147
                          `else
                            if(!1'b0) begin
                              $display("NOTE(SmartDispatcher.scala:147):    DEBUG-IDLE-FAST: First instruction is last in group (not branch/redirect), Group finished. -> IDLE"); // SmartDispatcher.scala:L147
                            end
                          `endif
                        `endif
                        isBusyReg <= 1'b0;
                        dispatchIndexReg <= 2'b00;
                      end else begin
                        dispatchIndexReg <= (io_fetchGroupIn_payload_startInstructionIndex + 2'b01);
                        `ifndef SYNTHESIS
                          `ifdef FORMAL
                            assert(1'b0); // SmartDispatcher.scala:L153
                          `else
                            if(!1'b0) begin
                              $display("NOTE(SmartDispatcher.scala:153):    DEBUG-IDLE-FAST: dispatchIndexReg set to %x + 1, FSM to DISPATCHING", dispatchIndexReg); // SmartDispatcher.scala:L153
                            end
                          `endif
                        `endif
                      end
                    end
                  end else begin
                    `ifndef SYNTHESIS
                      `ifdef FORMAL
                        assert(1'b0); // SmartDispatcher.scala:L158
                      `else
                        if(!1'b0) begin
                          $display("NOTE(SmartDispatcher.scala:158):  DISPATCHER-IDLE: First instruction (fast path) stalled. -> SEND_BRANCH"); // SmartDispatcher.scala:L158
                        end
                      `endif
                    `endif
                    `ifndef SYNTHESIS
                      `ifdef FORMAL
                        assert(1'b0); // SmartDispatcher.scala:L159
                      `else
                        if(!1'b0) begin
                          $display("NOTE(SmartDispatcher.scala:159):    DEBUG-IDLE-STALL: FSM to SEND_BRANCH"); // SmartDispatcher.scala:L159
                        end
                      `endif
                    `endif
                  end
                end else begin
                  `ifndef SYNTHESIS
                    `ifdef FORMAL
                      assert(1'b0); // SmartDispatcher.scala:L171
                    `else
                      if(!1'b0) begin
                        $display("NOTE(SmartDispatcher.scala:171):  DISPATCHER-IDLE: First instruction is Slow Path. PC=0x%x", _zz_io_fetchOutput_payload_pc); // SmartDispatcher.scala:L171
                      end
                    `endif
                  `endif
                  `ifndef SYNTHESIS
                    `ifdef FORMAL
                      assert(1'b0); // SmartDispatcher.scala:L185
                    `else
                      if(!1'b0) begin
                        $display("NOTE(SmartDispatcher.scala:185):  [notice] [33mDISPATCHER-IDLE: BPU Query sent for first instruction. -> WAITING_FOR_BPU[0m"); // SmartDispatcher.scala:L185
                      end
                    `endif
                  `endif
                end
              end
            end
          end
        end
        (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
          if(io_flush) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // SmartDispatcher.scala:L194
              `else
                if(!1'b0) begin
                  $display("NOTE(SmartDispatcher.scala:194):  [notice] [33mDISPATCHER: Flush received in DISPATCHING. -> DRAINING_BPU[0m"); // SmartDispatcher.scala:L194
                end
              `endif
            `endif
          end else begin
            if(isBusyReg) begin
              if(fetchGroupReg_fault) begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // SmartDispatcher.scala:L202
                  `else
                    if(!1'b0) begin
                      $display("NOTE(SmartDispatcher.scala:202):  DISPATCHER: Discarding faulted group PC=0x%x. -> IDLE", fetchGroupReg_pc); // SmartDispatcher.scala:L202
                    end
                  `endif
                `endif
                isBusyReg <= 1'b0;
                dispatchIndexReg <= 2'b00;
              end else begin
                if(when_SmartDispatcher_l206) begin
                  `ifndef SYNTHESIS
                    `ifdef FORMAL
                      assert(1'b0); // SmartDispatcher.scala:L207
                    `else
                      if(!1'b0) begin
                        $display("NOTE(SmartDispatcher.scala:207):  DISPATCHER: Complex Branch detected at PC=0x%x. -> QUERY_BPU", currentPcReg); // SmartDispatcher.scala:L207
                      end
                    `endif
                  `endif
                  `ifndef SYNTHESIS
                    `ifdef FORMAL
                      assert(1'b0); // SmartDispatcher.scala:L218
                    `else
                      if(!1'b0) begin
                        $display("NOTE(SmartDispatcher.scala:218):  DISPATCH-BURST: BPU Query sent for PC=0x%x. -> WAITING_FOR_BPU", currentPcReg); // SmartDispatcher.scala:L218
                      end
                    `endif
                  `endif
                end else begin
                  if(io_fetchOutput_ready) begin
                    `ifndef SYNTHESIS
                      `ifdef FORMAL
                        assert(1'b0); // SmartDispatcher.scala:L230
                      `else
                        if(!1'b0) begin
                          $display("NOTE(SmartDispatcher.scala:230):  DISPATCH-BURST: Fired PC=0x%x. isLast=%x, redirecting=%x", currentPcReg, isLastInstructionReg, currentPredecodeReg_isDirectJump); // SmartDispatcher.scala:L230
                        end
                      `endif
                    `endif
                    if(when_SmartDispatcher_l239) begin
                      `ifndef SYNTHESIS
                        `ifdef FORMAL
                          assert(1'b0); // SmartDispatcher.scala:L240
                        `else
                          if(!1'b0) begin
                            $display("NOTE(SmartDispatcher.scala:240):    DEBUG-DISPATCH-END: isLastInstruction=%x, redirecting=%x. Group finished. -> IDLE", isLastInstructionReg, currentPredecodeReg_isDirectJump); // SmartDispatcher.scala:L240
                          end
                        `endif
                      `endif
                      isBusyReg <= 1'b0;
                      dispatchIndexReg <= 2'b00;
                    end else begin
                      dispatchIndexReg <= (dispatchIndexReg + 2'b01);
                      `ifndef SYNTHESIS
                        `ifdef FORMAL
                          assert(1'b0); // SmartDispatcher.scala:L246
                        `else
                          if(!1'b0) begin
                            $display("NOTE(SmartDispatcher.scala:246):    DEBUG-DISPATCH-CONT: dispatchIndexReg set to %x + 1. Staying in DISPATCHING", dispatchIndexReg); // SmartDispatcher.scala:L246
                          end
                        `endif
                      `endif
                    end
                  end else begin
                    `ifndef SYNTHESIS
                      `ifdef FORMAL
                        assert(1'b0); // SmartDispatcher.scala:L250
                      `else
                        if(!1'b0) begin
                          $display("NOTE(SmartDispatcher.scala:250):  DISPATCH-BURST: Stalled for PC=0x%x", currentPcReg); // SmartDispatcher.scala:L250
                        end
                      `endif
                    `endif
                  end
                end
              end
            end else begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L254
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:254):  DISPATCHER-WARNING: isBusyReg is false but FSM is in DISPATCHING state. -> IDLE"); // SmartDispatcher.scala:L254
                  end
                `endif
              `endif
            end
          end
        end
        (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // SmartDispatcher.scala:L260
            `else
              if(!1'b0) begin
                $display("NOTE(SmartDispatcher.scala:260):  DISPATCH-WAIT-DEBUG: Current State (BEFORE flush check): io.flush=%x, io.bpuRsp.valid=%x, io.bpuRsp.payload.transactionId=%x, pendingTID=%x", io_flush, io_bpuRsp_valid, io_bpuRsp_payload_transactionId, pendingBpuQueryReg_bpuTransactionId); // SmartDispatcher.scala:L260
              end
            `endif
          `endif
          if(io_flush) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // SmartDispatcher.scala:L262
              `else
                if(!1'b0) begin
                  $display("NOTE(SmartDispatcher.scala:262):  [notice] [33mDISPATCHER: Flushing while WAITING_FOR_BPU. -> DRAINING_BPU[0m"); // SmartDispatcher.scala:L262
                end
              `endif
            `endif
          end else begin
            if(when_SmartDispatcher_l268) begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L269
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:269):  DISPATCH-WAIT: BPU Rsp mismatch because: valid=%x, transactionId=%x, pending=%x", io_bpuRsp_valid, io_bpuRsp_payload_transactionId, pendingBpuQueryReg_bpuTransactionId); // SmartDispatcher.scala:L269
                  end
                `endif
              `endif
            end
            if(when_SmartDispatcher_l273) begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L274
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:274):  DISPATCH-WAIT: Waiting BPU Rsp for PC=0x%x, TID=%x", pendingBpuQueryReg_pc, pendingBpuQueryReg_bpuTransactionId); // SmartDispatcher.scala:L274
                  end
                `endif
              `endif
            end
            if(when_SmartDispatcher_l279) begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L281
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:281):  [notice] [33mDISPATCH-WAIT: BPU Rsp Match! PC=0x%x, Taken=%x. -> SEND_BRANCH[0m", pendingBpuQueryReg_pc, io_bpuRsp_payload_isTaken); // SmartDispatcher.scala:L281
                  end
                `endif
              `endif
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L294
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:294):    DEBUG-OUTPUT-REG-UPDATED: outputReg.bpuPrediction.isTaken_ASSIGNED=%x, PC_ASSIGNED=%x", io_bpuRsp_payload_isTaken, pendingBpuQueryReg_pc); // SmartDispatcher.scala:L294
                  end
                `endif
              `endif
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L295
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:295):    DEBUG-OUTPUT-REG-UPDATED: outputReg.bpuPrediction.isTaken_REG_OUT=%x, PC_REG_OUT=%x", outputReg_bpuPrediction_isTaken, outputReg_pc); // SmartDispatcher.scala:L295
                  end
                `endif
              `endif
            end
          end
        end
        (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
          if(io_flush) begin
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // SmartDispatcher.scala:L304
              `else
                if(!1'b0) begin
                  $display("NOTE(SmartDispatcher.scala:304):  [notice] [33mDISPATCHER: Flush received in SEND_BRANCH. -> DRAINING_BPU[0m"); // SmartDispatcher.scala:L304
                end
              `endif
            `endif
          end else begin
            if(io_fetchOutput_fire) begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L312
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:312):  DISPATCH-SEND: Fired Branch/Stalled-FastPath PC=0x%x", outputReg_pc); // SmartDispatcher.scala:L312
                  end
                `endif
              `endif
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L313
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:313):    DEBUG-OUTPUT-FIRED: outputReg.bpuPrediction.isTaken=%x, PC=0x%x", outputReg_bpuPrediction_isTaken, outputReg_pc); // SmartDispatcher.scala:L313
                  end
                `endif
              `endif
              if(when_SmartDispatcher_l316) begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // SmartDispatcher.scala:L323
                  `else
                    if(!1'b0) begin
                      $display("NOTE(SmartDispatcher.scala:323):  DISPATCH-SEND: Soft redirect triggered to 0x%x", io_softRedirect_payload); // SmartDispatcher.scala:L323
                    end
                  `endif
                `endif
              end
              if(when_SmartDispatcher_l326) begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // SmartDispatcher.scala:L327
                  `else
                    if(!1'b0) begin
                      $display("NOTE(SmartDispatcher.scala:327):    DEBUG-SEND-END: isLastInstruction=%x, redirecting=%x. Group finished. -> IDLE", isLastInstructionReg, when_SmartDispatcher_l316); // SmartDispatcher.scala:L327
                    end
                  `endif
                `endif
                isBusyReg <= 1'b0;
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // SmartDispatcher.scala:L329
                  `else
                    if(!1'b0) begin
                      $display("NOTE(SmartDispatcher.scala:329):  DISPATCH-SEND: Group finished. -> IDLE"); // SmartDispatcher.scala:L329
                    end
                  `endif
                `endif
                dispatchIndexReg <= 2'b00;
              end else begin
                dispatchIndexReg <= (dispatchIndexReg + 2'b01);
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // SmartDispatcher.scala:L334
                  `else
                    if(!1'b0) begin
                      $display("NOTE(SmartDispatcher.scala:334):    DEBUG-SEND-CONT: dispatchIndexReg set to %x + 1. -> DISPATCHING", dispatchIndexReg); // SmartDispatcher.scala:L334
                    end
                  `endif
                `endif
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // SmartDispatcher.scala:L335
                  `else
                    if(!1'b0) begin
                      $display("NOTE(SmartDispatcher.scala:335):  DISPATCH-SEND: More instructions in group. -> DISPATCHING"); // SmartDispatcher.scala:L335
                    end
                  `endif
                `endif
              end
            end else begin
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L339
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:339):  DISPATCH-SEND: Stalled on output. PC=0x%x", outputReg_pc); // SmartDispatcher.scala:L339
                  end
                `endif
              `endif
              `ifndef SYNTHESIS
                `ifdef FORMAL
                  assert(1'b0); // SmartDispatcher.scala:L340
                `else
                  if(!1'b0) begin
                    $display("NOTE(SmartDispatcher.scala:340):    DEBUG-SEND-STALL: Stalled on output. PC=0x%x", outputReg_pc); // SmartDispatcher.scala:L340
                  end
                `endif
              `endif
            end
          end
        end
        (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // SmartDispatcher.scala:L346
            `else
              if(!1'b0) begin
                $display("NOTE(SmartDispatcher.scala:346):  DISPATCHER: Draining BPU requests. InFlight=%x", bpuInFlightCounterReg); // SmartDispatcher.scala:L346
              end
            `endif
          `endif
          if(when_SmartDispatcher_l347) begin
            isBusyReg <= 1'b0;
            dispatchIndexReg <= 2'b00;
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // SmartDispatcher.scala:L350
              `else
                if(!1'b0) begin
                  $display("NOTE(SmartDispatcher.scala:350):    DEBUG-ASSIGN: dispatchIndexReg assigned 0 from DRAINING_BPU"); // SmartDispatcher.scala:L350
                end
              `endif
            `endif
            `ifndef SYNTHESIS
              `ifdef FORMAL
                assert(1'b0); // SmartDispatcher.scala:L351
              `else
                if(!1'b0) begin
                  $display("NOTE(SmartDispatcher.scala:351):  DISPATCHER: BPU Draining complete. -> IDLE"); // SmartDispatcher.scala:L351
                end
              `endif
            `endif
          end
        end
        default : begin
        end
      endcase
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert(1'b0); // SmartDispatcher.scala:L365
        `else
          if(!1'b0) begin
            $display("NOTE(SmartDispatcher.scala:365):  DISPATCHER STATE: isBusyReg=%x, dispatchIndexReg=%x, fsmState=%s, bpuInFlight=%x", isBusyReg, dispatchIndexReg, fsm_stateReg_string, bpuInFlightCounterReg); // SmartDispatcher.scala:L365
          end
        `endif
      `endif
      if(io_fetchGroupIn_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // SmartDispatcher.scala:L368
          `else
            if(!1'b0) begin
              $display("NOTE(SmartDispatcher.scala:368):    -> EVENT: fetchGroupIn.fire"); // SmartDispatcher.scala:L368
            end
          `endif
        `endif
      end
      if(io_fetchOutput_fire) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // SmartDispatcher.scala:L369
          `else
            if(!1'b0) begin
              $display("NOTE(SmartDispatcher.scala:369):    -> EVENT: fetchOutput.fire"); // SmartDispatcher.scala:L369
            end
          `endif
        `endif
      end
      if(io_bpuQuery_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // SmartDispatcher.scala:L370
          `else
            if(!1'b0) begin
              $display("NOTE(SmartDispatcher.scala:370):    -> EVENT: bpuQuery.fire"); // SmartDispatcher.scala:L370
            end
          `endif
        `endif
      end
      if(io_bpuRsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // SmartDispatcher.scala:L371
          `else
            if(!1'b0) begin
              $display("NOTE(SmartDispatcher.scala:371):    -> EVENT: bpuRsp.fire"); // SmartDispatcher.scala:L371
            end
          `endif
        `endif
      end
      if(io_softRedirect_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // SmartDispatcher.scala:L372
          `else
            if(!1'b0) begin
              $display("NOTE(SmartDispatcher.scala:372):    -> EVENT: softRedirect.valid"); // SmartDispatcher.scala:L372
            end
          `endif
        `endif
      end
      if(io_flush) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // SmartDispatcher.scala:L373
          `else
            if(!1'b0) begin
              $display("NOTE(SmartDispatcher.scala:373):    -> EVENT: FLUSH asserted"); // SmartDispatcher.scala:L373
            end
          `endif
        `endif
      end
    end
  end

  always @(posedge clk) begin
    if(io_flush) begin
      fetchGroupReg_pc <= 32'h0;
      fetchGroupReg_instructions_0 <= 32'h0;
      fetchGroupReg_instructions_1 <= 32'h0;
      fetchGroupReg_instructions_2 <= 32'h0;
      fetchGroupReg_instructions_3 <= 32'h0;
      fetchGroupReg_predecodeInfos_0_isBranch <= 1'b0;
      fetchGroupReg_predecodeInfos_0_isJump <= 1'b0;
      fetchGroupReg_predecodeInfos_0_isDirectJump <= 1'b0;
      fetchGroupReg_predecodeInfos_0_jumpOffset <= 32'h0;
      fetchGroupReg_predecodeInfos_0_isIdle <= 1'b0;
      fetchGroupReg_predecodeInfos_1_isBranch <= 1'b0;
      fetchGroupReg_predecodeInfos_1_isJump <= 1'b0;
      fetchGroupReg_predecodeInfos_1_isDirectJump <= 1'b0;
      fetchGroupReg_predecodeInfos_1_jumpOffset <= 32'h0;
      fetchGroupReg_predecodeInfos_1_isIdle <= 1'b0;
      fetchGroupReg_predecodeInfos_2_isBranch <= 1'b0;
      fetchGroupReg_predecodeInfos_2_isJump <= 1'b0;
      fetchGroupReg_predecodeInfos_2_isDirectJump <= 1'b0;
      fetchGroupReg_predecodeInfos_2_jumpOffset <= 32'h0;
      fetchGroupReg_predecodeInfos_2_isIdle <= 1'b0;
      fetchGroupReg_predecodeInfos_3_isBranch <= 1'b0;
      fetchGroupReg_predecodeInfos_3_isJump <= 1'b0;
      fetchGroupReg_predecodeInfos_3_isDirectJump <= 1'b0;
      fetchGroupReg_predecodeInfos_3_jumpOffset <= 32'h0;
      fetchGroupReg_predecodeInfos_3_isIdle <= 1'b0;
      fetchGroupReg_branchMask <= 4'b0000;
      fetchGroupReg_fault <= 1'b0;
      fetchGroupReg_numValidInstructions <= 3'b000;
      fetchGroupReg_startInstructionIndex <= 2'b00;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (fsm_stateReg[fsm_1_IDLE_OH_ID]) : begin
        if(!io_flush) begin
          if(io_fetchGroupIn_fire) begin
            fetchGroupReg_pc <= io_fetchGroupIn_payload_pc;
            fetchGroupReg_instructions_0 <= io_fetchGroupIn_payload_instructions_0;
            fetchGroupReg_instructions_1 <= io_fetchGroupIn_payload_instructions_1;
            fetchGroupReg_instructions_2 <= io_fetchGroupIn_payload_instructions_2;
            fetchGroupReg_instructions_3 <= io_fetchGroupIn_payload_instructions_3;
            fetchGroupReg_predecodeInfos_0_isBranch <= io_fetchGroupIn_payload_predecodeInfos_0_isBranch;
            fetchGroupReg_predecodeInfos_0_isJump <= io_fetchGroupIn_payload_predecodeInfos_0_isJump;
            fetchGroupReg_predecodeInfos_0_isDirectJump <= io_fetchGroupIn_payload_predecodeInfos_0_isDirectJump;
            fetchGroupReg_predecodeInfos_0_jumpOffset <= io_fetchGroupIn_payload_predecodeInfos_0_jumpOffset;
            fetchGroupReg_predecodeInfos_0_isIdle <= io_fetchGroupIn_payload_predecodeInfos_0_isIdle;
            fetchGroupReg_predecodeInfos_1_isBranch <= io_fetchGroupIn_payload_predecodeInfos_1_isBranch;
            fetchGroupReg_predecodeInfos_1_isJump <= io_fetchGroupIn_payload_predecodeInfos_1_isJump;
            fetchGroupReg_predecodeInfos_1_isDirectJump <= io_fetchGroupIn_payload_predecodeInfos_1_isDirectJump;
            fetchGroupReg_predecodeInfos_1_jumpOffset <= io_fetchGroupIn_payload_predecodeInfos_1_jumpOffset;
            fetchGroupReg_predecodeInfos_1_isIdle <= io_fetchGroupIn_payload_predecodeInfos_1_isIdle;
            fetchGroupReg_predecodeInfos_2_isBranch <= io_fetchGroupIn_payload_predecodeInfos_2_isBranch;
            fetchGroupReg_predecodeInfos_2_isJump <= io_fetchGroupIn_payload_predecodeInfos_2_isJump;
            fetchGroupReg_predecodeInfos_2_isDirectJump <= io_fetchGroupIn_payload_predecodeInfos_2_isDirectJump;
            fetchGroupReg_predecodeInfos_2_jumpOffset <= io_fetchGroupIn_payload_predecodeInfos_2_jumpOffset;
            fetchGroupReg_predecodeInfos_2_isIdle <= io_fetchGroupIn_payload_predecodeInfos_2_isIdle;
            fetchGroupReg_predecodeInfos_3_isBranch <= io_fetchGroupIn_payload_predecodeInfos_3_isBranch;
            fetchGroupReg_predecodeInfos_3_isJump <= io_fetchGroupIn_payload_predecodeInfos_3_isJump;
            fetchGroupReg_predecodeInfos_3_isDirectJump <= io_fetchGroupIn_payload_predecodeInfos_3_isDirectJump;
            fetchGroupReg_predecodeInfos_3_jumpOffset <= io_fetchGroupIn_payload_predecodeInfos_3_jumpOffset;
            fetchGroupReg_predecodeInfos_3_isIdle <= io_fetchGroupIn_payload_predecodeInfos_3_isIdle;
            fetchGroupReg_branchMask <= io_fetchGroupIn_payload_branchMask;
            fetchGroupReg_fault <= io_fetchGroupIn_payload_fault;
            fetchGroupReg_numValidInstructions <= io_fetchGroupIn_payload_numValidInstructions;
            fetchGroupReg_startInstructionIndex <= io_fetchGroupIn_payload_startInstructionIndex;
            if(!when_SmartDispatcher_l108) begin
              if(when_SmartDispatcher_l123) begin
                if(!io_fetchOutput_ready) begin
                  outputReg_pc <= _zz_io_fetchOutput_payload_pc;
                  outputReg_instruction <= _zz_io_fetchOutput_payload_instruction;
                  outputReg_predecode_isBranch <= _zz_io_fetchOutput_payload_predecode_isBranch;
                  outputReg_predecode_isJump <= _zz_io_fetchOutput_payload_predecode_isJump;
                  outputReg_predecode_isDirectJump <= _zz_io_fetchOutput_payload_predecode_isDirectJump;
                  outputReg_predecode_jumpOffset <= _zz_io_fetchOutput_payload_predecode_jumpOffset;
                  outputReg_predecode_isIdle <= _zz_io_fetchOutput_payload_predecode_isIdle;
                  outputReg_bpuPrediction_isTaken <= 1'b0;
                  outputReg_bpuPrediction_target <= 32'h0;
                  outputReg_bpuPrediction_wasPredicted <= 1'b0;
                end
              end else begin
                pendingBpuQueryReg_pc <= _zz_io_fetchOutput_payload_pc;
                pendingBpuQueryReg_instruction <= _zz_io_fetchOutput_payload_instruction;
                pendingBpuQueryReg_predecodeInfo_isBranch <= _zz_io_fetchOutput_payload_predecode_isBranch;
                pendingBpuQueryReg_predecodeInfo_isJump <= _zz_io_fetchOutput_payload_predecode_isJump;
                pendingBpuQueryReg_predecodeInfo_isDirectJump <= _zz_io_fetchOutput_payload_predecode_isDirectJump;
                pendingBpuQueryReg_predecodeInfo_jumpOffset <= _zz_io_fetchOutput_payload_predecode_jumpOffset;
                pendingBpuQueryReg_predecodeInfo_isIdle <= _zz_io_fetchOutput_payload_predecode_isIdle;
                pendingBpuQueryReg_bpuTransactionId <= bpuTransIdCounterReg;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_DISPATCHING_OH_ID]) : begin
        if(!io_flush) begin
          if(isBusyReg) begin
            if(!fetchGroupReg_fault) begin
              if(when_SmartDispatcher_l206) begin
                pendingBpuQueryReg_pc <= currentPcReg;
                pendingBpuQueryReg_instruction <= currentInstructionReg;
                pendingBpuQueryReg_predecodeInfo_isBranch <= currentPredecodeReg_isBranch;
                pendingBpuQueryReg_predecodeInfo_isJump <= currentPredecodeReg_isJump;
                pendingBpuQueryReg_predecodeInfo_isDirectJump <= currentPredecodeReg_isDirectJump;
                pendingBpuQueryReg_predecodeInfo_jumpOffset <= currentPredecodeReg_jumpOffset;
                pendingBpuQueryReg_predecodeInfo_isIdle <= currentPredecodeReg_isIdle;
                pendingBpuQueryReg_bpuTransactionId <= bpuTransIdCounterReg;
              end
            end
          end
        end
      end
      (fsm_stateReg[fsm_1_WAITING_FOR_BPU_OH_ID]) : begin
        if(!io_flush) begin
          if(when_SmartDispatcher_l279) begin
            outputReg_pc <= pendingBpuQueryReg_pc;
            outputReg_instruction <= pendingBpuQueryReg_instruction;
            outputReg_predecode_isBranch <= pendingBpuQueryReg_predecodeInfo_isBranch;
            outputReg_predecode_isJump <= pendingBpuQueryReg_predecodeInfo_isJump;
            outputReg_predecode_isDirectJump <= pendingBpuQueryReg_predecodeInfo_isDirectJump;
            outputReg_predecode_jumpOffset <= pendingBpuQueryReg_predecodeInfo_jumpOffset;
            outputReg_predecode_isIdle <= pendingBpuQueryReg_predecodeInfo_isIdle;
            outputReg_bpuPrediction_wasPredicted <= 1'b1;
            outputReg_bpuPrediction_isTaken <= io_bpuRsp_payload_isTaken;
            outputReg_bpuPrediction_target <= io_bpuRsp_payload_target;
          end
        end
      end
      (fsm_stateReg[fsm_1_SEND_BRANCH_OH_ID]) : begin
      end
      (fsm_stateReg[fsm_1_DRAINING_BPU_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end


endmodule

//OneShot_12 replaced by OneShot

module StreamArbiter_7 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [3:0]    io_inputs_0_payload_robPtr,
  input  wire [5:0]    io_inputs_0_payload_pdest,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire          io_inputs_0_payload_isIO,
  input  wire [1:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_hasEarlyException,
  input  wire [7:0]    io_inputs_0_payload_earlyExceptionCode,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [3:0]    io_output_payload_robPtr,
  output wire [5:0]    io_output_payload_pdest,
  output wire [31:0]   io_output_payload_address,
  output wire          io_output_payload_isIO,
  output wire [1:0]    io_output_payload_size,
  output wire          io_output_payload_hasEarlyException,
  output wire [7:0]    io_output_payload_earlyExceptionCode,
  output wire [0:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;
  wire                io_output_fire;
  wire       [1:0]    _zz_io_output_payload_size;
  `ifndef SYNTHESIS
  reg [7:0] io_inputs_0_payload_size_string;
  reg [7:0] io_output_payload_size_string;
  reg [7:0] _zz_io_output_payload_size_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_size)
      MemAccessSize_B : io_inputs_0_payload_size_string = "B";
      MemAccessSize_H : io_inputs_0_payload_size_string = "H";
      MemAccessSize_W : io_inputs_0_payload_size_string = "W";
      MemAccessSize_D : io_inputs_0_payload_size_string = "D";
      default : io_inputs_0_payload_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_output_payload_size)
      MemAccessSize_B : io_output_payload_size_string = "B";
      MemAccessSize_H : io_output_payload_size_string = "H";
      MemAccessSize_W : io_output_payload_size_string = "W";
      MemAccessSize_D : io_output_payload_size_string = "D";
      default : io_output_payload_size_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_size)
      MemAccessSize_B : _zz_io_output_payload_size_string = "B";
      MemAccessSize_H : _zz_io_output_payload_size_string = "H";
      MemAccessSize_W : _zz_io_output_payload_size_string = "W";
      MemAccessSize_D : _zz_io_output_payload_size_string = "D";
      default : _zz_io_output_payload_size_string = "?";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign _zz_io_output_payload_size = io_inputs_0_payload_size;
  assign io_output_payload_robPtr = io_inputs_0_payload_robPtr;
  assign io_output_payload_pdest = io_inputs_0_payload_pdest;
  assign io_output_payload_address = io_inputs_0_payload_address;
  assign io_output_payload_isIO = io_inputs_0_payload_isIO;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_hasEarlyException = io_inputs_0_payload_hasEarlyException;
  assign io_output_payload_earlyExceptionCode = io_inputs_0_payload_earlyExceptionCode;
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk) begin
    if(reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

//OneShot_11 replaced by OneShot

module StreamDemux (
  input  wire [0:0]    io_select,
  input  wire          io_input_valid,
  output reg           io_input_ready,
  input  wire [2:0]    io_input_payload_qPtr,
  input  wire [31:0]   io_input_payload_address,
  input  wire          io_input_payload_alignException,
  input  wire [1:0]    io_input_payload_accessSize,
  input  wire [3:0]    io_input_payload_storeMask,
  input  wire [5:0]    io_input_payload_basePhysReg,
  input  wire [31:0]   io_input_payload_immediate,
  input  wire          io_input_payload_usePc,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [3:0]    io_input_payload_robPtr,
  input  wire          io_input_payload_isLoad,
  input  wire          io_input_payload_isStore,
  input  wire [5:0]    io_input_payload_physDst,
  input  wire [31:0]   io_input_payload_storeData,
  input  wire          io_input_payload_isFlush,
  input  wire          io_input_payload_isIO,
  output reg           io_outputs_0_valid,
  input  wire          io_outputs_0_ready,
  output wire [2:0]    io_outputs_0_payload_qPtr,
  output wire [31:0]   io_outputs_0_payload_address,
  output wire          io_outputs_0_payload_alignException,
  output wire [1:0]    io_outputs_0_payload_accessSize,
  output wire [3:0]    io_outputs_0_payload_storeMask,
  output wire [5:0]    io_outputs_0_payload_basePhysReg,
  output wire [31:0]   io_outputs_0_payload_immediate,
  output wire          io_outputs_0_payload_usePc,
  output wire [31:0]   io_outputs_0_payload_pc,
  output wire [3:0]    io_outputs_0_payload_robPtr,
  output wire          io_outputs_0_payload_isLoad,
  output wire          io_outputs_0_payload_isStore,
  output wire [5:0]    io_outputs_0_payload_physDst,
  output wire [31:0]   io_outputs_0_payload_storeData,
  output wire          io_outputs_0_payload_isFlush,
  output wire          io_outputs_0_payload_isIO,
  output reg           io_outputs_1_valid,
  input  wire          io_outputs_1_ready,
  output wire [2:0]    io_outputs_1_payload_qPtr,
  output wire [31:0]   io_outputs_1_payload_address,
  output wire          io_outputs_1_payload_alignException,
  output wire [1:0]    io_outputs_1_payload_accessSize,
  output wire [3:0]    io_outputs_1_payload_storeMask,
  output wire [5:0]    io_outputs_1_payload_basePhysReg,
  output wire [31:0]   io_outputs_1_payload_immediate,
  output wire          io_outputs_1_payload_usePc,
  output wire [31:0]   io_outputs_1_payload_pc,
  output wire [3:0]    io_outputs_1_payload_robPtr,
  output wire          io_outputs_1_payload_isLoad,
  output wire          io_outputs_1_payload_isStore,
  output wire [5:0]    io_outputs_1_payload_physDst,
  output wire [31:0]   io_outputs_1_payload_storeData,
  output wire          io_outputs_1_payload_isFlush,
  output wire          io_outputs_1_payload_isIO
);
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;

  wire                when_Stream_l1168;
  wire                when_Stream_l1168_1;
  `ifndef SYNTHESIS
  reg [7:0] io_input_payload_accessSize_string;
  reg [7:0] io_outputs_0_payload_accessSize_string;
  reg [7:0] io_outputs_1_payload_accessSize_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_accessSize)
      MemAccessSize_B : io_input_payload_accessSize_string = "B";
      MemAccessSize_H : io_input_payload_accessSize_string = "H";
      MemAccessSize_W : io_input_payload_accessSize_string = "W";
      MemAccessSize_D : io_input_payload_accessSize_string = "D";
      default : io_input_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_payload_accessSize)
      MemAccessSize_B : io_outputs_0_payload_accessSize_string = "B";
      MemAccessSize_H : io_outputs_0_payload_accessSize_string = "H";
      MemAccessSize_W : io_outputs_0_payload_accessSize_string = "W";
      MemAccessSize_D : io_outputs_0_payload_accessSize_string = "D";
      default : io_outputs_0_payload_accessSize_string = "?";
    endcase
  end
  always @(*) begin
    case(io_outputs_1_payload_accessSize)
      MemAccessSize_B : io_outputs_1_payload_accessSize_string = "B";
      MemAccessSize_H : io_outputs_1_payload_accessSize_string = "H";
      MemAccessSize_W : io_outputs_1_payload_accessSize_string = "W";
      MemAccessSize_D : io_outputs_1_payload_accessSize_string = "D";
      default : io_outputs_1_payload_accessSize_string = "?";
    endcase
  end
  `endif

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l1168) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l1168_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_qPtr = io_input_payload_qPtr;
  assign io_outputs_0_payload_address = io_input_payload_address;
  assign io_outputs_0_payload_alignException = io_input_payload_alignException;
  assign io_outputs_0_payload_accessSize = io_input_payload_accessSize;
  assign io_outputs_0_payload_storeMask = io_input_payload_storeMask;
  assign io_outputs_0_payload_basePhysReg = io_input_payload_basePhysReg;
  assign io_outputs_0_payload_immediate = io_input_payload_immediate;
  assign io_outputs_0_payload_usePc = io_input_payload_usePc;
  assign io_outputs_0_payload_pc = io_input_payload_pc;
  assign io_outputs_0_payload_robPtr = io_input_payload_robPtr;
  assign io_outputs_0_payload_isLoad = io_input_payload_isLoad;
  assign io_outputs_0_payload_isStore = io_input_payload_isStore;
  assign io_outputs_0_payload_physDst = io_input_payload_physDst;
  assign io_outputs_0_payload_storeData = io_input_payload_storeData;
  assign io_outputs_0_payload_isFlush = io_input_payload_isFlush;
  assign io_outputs_0_payload_isIO = io_input_payload_isIO;
  assign when_Stream_l1168 = (1'b0 != io_select);
  always @(*) begin
    if(when_Stream_l1168) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_qPtr = io_input_payload_qPtr;
  assign io_outputs_1_payload_address = io_input_payload_address;
  assign io_outputs_1_payload_alignException = io_input_payload_alignException;
  assign io_outputs_1_payload_accessSize = io_input_payload_accessSize;
  assign io_outputs_1_payload_storeMask = io_input_payload_storeMask;
  assign io_outputs_1_payload_basePhysReg = io_input_payload_basePhysReg;
  assign io_outputs_1_payload_immediate = io_input_payload_immediate;
  assign io_outputs_1_payload_usePc = io_input_payload_usePc;
  assign io_outputs_1_payload_pc = io_input_payload_pc;
  assign io_outputs_1_payload_robPtr = io_input_payload_robPtr;
  assign io_outputs_1_payload_isLoad = io_input_payload_isLoad;
  assign io_outputs_1_payload_isStore = io_input_payload_isStore;
  assign io_outputs_1_payload_physDst = io_input_payload_physDst;
  assign io_outputs_1_payload_storeData = io_input_payload_storeData;
  assign io_outputs_1_payload_isFlush = io_input_payload_isFlush;
  assign io_outputs_1_payload_isIO = io_input_payload_isIO;
  assign when_Stream_l1168_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Stream_l1168_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

//OneShot_10 replaced by OneShot

//OneShot_9 replaced by OneShot

//OneShot_8 replaced by OneShot

module FrequencyDivider (
  output wire          io_tick,
  input  wire          clk,
  input  wire          reset
);

  reg        [26:0]   counter;

  assign io_tick = (counter == 27'h5f5e0ff);
  always @(posedge clk) begin
    if(reset) begin
      counter <= 27'h0;
    end else begin
      if(io_tick) begin
        counter <= 27'h0;
      end else begin
        counter <= (counter + 27'h0000001);
      end
    end
  end


endmodule

//OneShot_7 replaced by OneShot

module IssueQueueComponent_3 (
  input  wire          io_allocateIn_valid,
  output wire          io_allocateIn_ready,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_pc,
  input  wire          io_allocateIn_payload_uop_decoded_isValid,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_uopCode,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_exeUnit,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_isa,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archDest_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archDest_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_writeArchDestEn,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archSrc1_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archSrc1_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_useArchSrc1,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archSrc2_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archSrc2_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_useArchSrc2,
  input  wire          io_allocateIn_payload_uop_decoded_usePcForAddr,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_imm,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_immUsage,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isSub,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isAdd,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isSigned,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_aluCtrl_logicOp,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isRight,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_memCtrl_size,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isStore,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_memCtrl_atomicOp,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isFence,
  input  wire [7:0]    io_allocateIn_payload_uop_decoded_memCtrl_fenceMode,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_branchCtrl_condition,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isJump,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isLink,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_opType,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond,
  input  wire [13:0]   io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isWrite,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isRead,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isExchange,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc,
  input  wire [19:0]   io_allocateIn_payload_uop_decoded_sysCtrl_sysCode,
  input  wire          io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn,
  input  wire          io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_decodeExceptionCode,
  input  wire          io_allocateIn_payload_uop_decoded_hasDecodeException,
  input  wire          io_allocateIn_payload_uop_decoded_isMicrocode,
  input  wire [7:0]    io_allocateIn_payload_uop_decoded_microcodeEntry,
  input  wire          io_allocateIn_payload_uop_decoded_isSerializing,
  input  wire          io_allocateIn_payload_uop_decoded_isBranchOrJump,
  input  wire          io_allocateIn_payload_uop_decoded_branchPrediction_isTaken,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_branchPrediction_target,
  input  wire          io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physSrc1_idx,
  input  wire          io_allocateIn_payload_uop_rename_physSrc1IsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physSrc2_idx,
  input  wire          io_allocateIn_payload_uop_rename_physSrc2IsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physDest_idx,
  input  wire          io_allocateIn_payload_uop_rename_physDestIsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_oldPhysDest_idx,
  input  wire          io_allocateIn_payload_uop_rename_oldPhysDestIsFpr,
  input  wire          io_allocateIn_payload_uop_rename_allocatesPhysDest,
  input  wire          io_allocateIn_payload_uop_rename_writesToPhysReg,
  input  wire [3:0]    io_allocateIn_payload_uop_robPtr,
  input  wire [15:0]   io_allocateIn_payload_uop_uniqueId,
  input  wire          io_allocateIn_payload_uop_dispatched,
  input  wire          io_allocateIn_payload_uop_executed,
  input  wire          io_allocateIn_payload_uop_hasException,
  input  wire [7:0]    io_allocateIn_payload_uop_exceptionCode,
  input  wire          io_allocateIn_payload_src1InitialReady,
  input  wire          io_allocateIn_payload_src2InitialReady,
  output wire          io_issueOut_valid,
  input  wire          io_issueOut_ready,
  output wire [3:0]    io_issueOut_payload_robPtr,
  output wire [5:0]    io_issueOut_payload_physDest_idx,
  output wire          io_issueOut_payload_physDestIsFpr,
  output wire          io_issueOut_payload_writesToPhysReg,
  output wire          io_issueOut_payload_useSrc1,
  output wire [31:0]   io_issueOut_payload_src1Data,
  output wire [5:0]    io_issueOut_payload_src1Tag,
  output wire          io_issueOut_payload_src1Ready,
  output wire          io_issueOut_payload_src1IsFpr,
  output wire          io_issueOut_payload_useSrc2,
  output wire [31:0]   io_issueOut_payload_src2Data,
  output wire [5:0]    io_issueOut_payload_src2Tag,
  output wire          io_issueOut_payload_src2Ready,
  output wire          io_issueOut_payload_src2IsFpr,
  output wire [1:0]    io_issueOut_payload_memCtrl_size,
  output wire          io_issueOut_payload_memCtrl_isSignedLoad,
  output wire          io_issueOut_payload_memCtrl_isStore,
  output wire          io_issueOut_payload_memCtrl_isLoadLinked,
  output wire          io_issueOut_payload_memCtrl_isStoreCond,
  output wire [4:0]    io_issueOut_payload_memCtrl_atomicOp,
  output wire          io_issueOut_payload_memCtrl_isFence,
  output wire [7:0]    io_issueOut_payload_memCtrl_fenceMode,
  output wire          io_issueOut_payload_memCtrl_isCacheOp,
  output wire [4:0]    io_issueOut_payload_memCtrl_cacheOpType,
  output wire          io_issueOut_payload_memCtrl_isPrefetch,
  output wire [31:0]   io_issueOut_payload_imm,
  output wire          io_issueOut_payload_usePc,
  output wire [31:0]   io_issueOut_payload_pcData,
  input  wire          io_wakeupIn_0_valid,
  input  wire [5:0]    io_wakeupIn_0_payload_physRegIdx,
  input  wire          io_wakeupIn_1_valid,
  input  wire [5:0]    io_wakeupIn_1_payload_physRegIdx,
  input  wire          io_wakeupIn_2_valid,
  input  wire [5:0]    io_wakeupIn_2_payload_physRegIdx,
  input  wire          io_wakeupIn_3_valid,
  input  wire [5:0]    io_wakeupIn_3_payload_physRegIdx,
  input  wire          io_wakeupIn_4_valid,
  input  wire [5:0]    io_wakeupIn_4_payload_physRegIdx,
  input  wire          io_flush,
  input  wire          clk,
  input  wire          reset
);
  localparam BaseUopCode_NOP = 5'd0;
  localparam BaseUopCode_ILLEGAL = 5'd1;
  localparam BaseUopCode_ALU = 5'd2;
  localparam BaseUopCode_SHIFT = 5'd3;
  localparam BaseUopCode_MUL = 5'd4;
  localparam BaseUopCode_DIV = 5'd5;
  localparam BaseUopCode_LOAD = 5'd6;
  localparam BaseUopCode_STORE = 5'd7;
  localparam BaseUopCode_ATOMIC = 5'd8;
  localparam BaseUopCode_MEM_BARRIER = 5'd9;
  localparam BaseUopCode_PREFETCH = 5'd10;
  localparam BaseUopCode_BRANCH = 5'd11;
  localparam BaseUopCode_JUMP_REG = 5'd12;
  localparam BaseUopCode_JUMP_IMM = 5'd13;
  localparam BaseUopCode_SYSTEM_OP = 5'd14;
  localparam BaseUopCode_CSR_ACCESS = 5'd15;
  localparam BaseUopCode_FPU_ALU = 5'd16;
  localparam BaseUopCode_FPU_CVT = 5'd17;
  localparam BaseUopCode_FPU_CMP = 5'd18;
  localparam BaseUopCode_FPU_SEL = 5'd19;
  localparam BaseUopCode_LA_BITMANIP = 5'd20;
  localparam BaseUopCode_LA_CACOP = 5'd21;
  localparam BaseUopCode_LA_TLB = 5'd22;
  localparam BaseUopCode_IDLE = 5'd23;
  localparam ExeUnitType_NONE = 4'd0;
  localparam ExeUnitType_ALU_INT = 4'd1;
  localparam ExeUnitType_MUL_INT = 4'd2;
  localparam ExeUnitType_DIV_INT = 4'd3;
  localparam ExeUnitType_MEM = 4'd4;
  localparam ExeUnitType_BRU = 4'd5;
  localparam ExeUnitType_CSR = 4'd6;
  localparam ExeUnitType_FPU_ADD_MUL_CVT_CMP = 4'd7;
  localparam ExeUnitType_FPU_DIV_SQRT = 4'd8;
  localparam IsaType_UNKNOWN = 2'd0;
  localparam IsaType_DEMO = 2'd1;
  localparam IsaType_RISCV = 2'd2;
  localparam IsaType_LOONGARCH = 2'd3;
  localparam ArchRegType_GPR = 2'd0;
  localparam ArchRegType_FPR = 2'd1;
  localparam ArchRegType_CSR = 2'd2;
  localparam ArchRegType_LA_CF = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;
  localparam BranchCondition_NUL = 5'd0;
  localparam BranchCondition_EQ = 5'd1;
  localparam BranchCondition_NE = 5'd2;
  localparam BranchCondition_LT = 5'd3;
  localparam BranchCondition_GE = 5'd4;
  localparam BranchCondition_LTU = 5'd5;
  localparam BranchCondition_GEU = 5'd6;
  localparam BranchCondition_EQZ = 5'd7;
  localparam BranchCondition_NEZ = 5'd8;
  localparam BranchCondition_LTZ = 5'd9;
  localparam BranchCondition_GEZ = 5'd10;
  localparam BranchCondition_GTZ = 5'd11;
  localparam BranchCondition_LEZ = 5'd12;
  localparam BranchCondition_F_EQ = 5'd13;
  localparam BranchCondition_F_NE = 5'd14;
  localparam BranchCondition_F_LT = 5'd15;
  localparam BranchCondition_F_LE = 5'd16;
  localparam BranchCondition_F_UN = 5'd17;
  localparam BranchCondition_LA_CF_TRUE = 5'd18;
  localparam BranchCondition_LA_CF_FALSE = 5'd19;
  localparam DecodeExCode_INVALID = 2'd0;
  localparam DecodeExCode_FETCH_ERROR = 2'd1;
  localparam DecodeExCode_DECODE_ERROR = 2'd2;
  localparam DecodeExCode_OK = 2'd3;

  wire       [3:0]    _zz_issueRequestMask_ohFirst_masked;
  reg        [1:0]    _zz__zz_io_issueOut_payload_memCtrl_size;
  reg        [3:0]    _zz_io_issueOut_payload_robPtr;
  reg        [5:0]    _zz_io_issueOut_payload_physDest_idx;
  reg                 _zz_io_issueOut_payload_physDestIsFpr;
  reg                 _zz_io_issueOut_payload_writesToPhysReg;
  reg                 _zz_io_issueOut_payload_useSrc1;
  reg        [31:0]   _zz_io_issueOut_payload_src1Data;
  reg        [5:0]    _zz_io_issueOut_payload_src1Tag;
  reg                 _zz_io_issueOut_payload_src1Ready;
  reg                 _zz_io_issueOut_payload_src1IsFpr;
  reg                 _zz_io_issueOut_payload_useSrc2;
  reg        [31:0]   _zz_io_issueOut_payload_src2Data;
  reg        [5:0]    _zz_io_issueOut_payload_src2Tag;
  reg                 _zz_io_issueOut_payload_src2Ready;
  reg                 _zz_io_issueOut_payload_src2IsFpr;
  reg                 _zz_io_issueOut_payload_memCtrl_isSignedLoad;
  reg                 _zz_io_issueOut_payload_memCtrl_isStore;
  reg                 _zz_io_issueOut_payload_memCtrl_isLoadLinked;
  reg                 _zz_io_issueOut_payload_memCtrl_isStoreCond;
  reg        [4:0]    _zz_io_issueOut_payload_memCtrl_atomicOp;
  reg                 _zz_io_issueOut_payload_memCtrl_isFence;
  reg        [7:0]    _zz_io_issueOut_payload_memCtrl_fenceMode;
  reg                 _zz_io_issueOut_payload_memCtrl_isCacheOp;
  reg        [4:0]    _zz_io_issueOut_payload_memCtrl_cacheOpType;
  reg                 _zz_io_issueOut_payload_memCtrl_isPrefetch;
  reg        [31:0]   _zz_io_issueOut_payload_imm;
  reg                 _zz_io_issueOut_payload_usePc;
  reg        [31:0]   _zz_io_issueOut_payload_pcData;
  wire       [3:0]    _zz_allocationMask_1;
  reg        [2:0]    _zz_currentValidCount_8;
  wire       [2:0]    _zz_currentValidCount_9;
  reg        [2:0]    _zz_currentValidCount_10;
  wire       [2:0]    _zz_currentValidCount_11;
  wire       [0:0]    _zz_currentValidCount_12;
  reg        [3:0]    entries_0_robPtr;
  reg        [5:0]    entries_0_physDest_idx;
  reg                 entries_0_physDestIsFpr;
  reg                 entries_0_writesToPhysReg;
  reg                 entries_0_useSrc1;
  reg        [31:0]   entries_0_src1Data;
  reg        [5:0]    entries_0_src1Tag;
  reg                 entries_0_src1Ready;
  reg                 entries_0_src1IsFpr;
  reg                 entries_0_useSrc2;
  reg        [31:0]   entries_0_src2Data;
  reg        [5:0]    entries_0_src2Tag;
  reg                 entries_0_src2Ready;
  reg                 entries_0_src2IsFpr;
  reg        [1:0]    entries_0_memCtrl_size;
  reg                 entries_0_memCtrl_isSignedLoad;
  reg                 entries_0_memCtrl_isStore;
  reg                 entries_0_memCtrl_isLoadLinked;
  reg                 entries_0_memCtrl_isStoreCond;
  reg        [4:0]    entries_0_memCtrl_atomicOp;
  reg                 entries_0_memCtrl_isFence;
  reg        [7:0]    entries_0_memCtrl_fenceMode;
  reg                 entries_0_memCtrl_isCacheOp;
  reg        [4:0]    entries_0_memCtrl_cacheOpType;
  reg                 entries_0_memCtrl_isPrefetch;
  reg        [31:0]   entries_0_imm;
  reg                 entries_0_usePc;
  reg        [31:0]   entries_0_pcData;
  reg        [3:0]    entries_1_robPtr;
  reg        [5:0]    entries_1_physDest_idx;
  reg                 entries_1_physDestIsFpr;
  reg                 entries_1_writesToPhysReg;
  reg                 entries_1_useSrc1;
  reg        [31:0]   entries_1_src1Data;
  reg        [5:0]    entries_1_src1Tag;
  reg                 entries_1_src1Ready;
  reg                 entries_1_src1IsFpr;
  reg                 entries_1_useSrc2;
  reg        [31:0]   entries_1_src2Data;
  reg        [5:0]    entries_1_src2Tag;
  reg                 entries_1_src2Ready;
  reg                 entries_1_src2IsFpr;
  reg        [1:0]    entries_1_memCtrl_size;
  reg                 entries_1_memCtrl_isSignedLoad;
  reg                 entries_1_memCtrl_isStore;
  reg                 entries_1_memCtrl_isLoadLinked;
  reg                 entries_1_memCtrl_isStoreCond;
  reg        [4:0]    entries_1_memCtrl_atomicOp;
  reg                 entries_1_memCtrl_isFence;
  reg        [7:0]    entries_1_memCtrl_fenceMode;
  reg                 entries_1_memCtrl_isCacheOp;
  reg        [4:0]    entries_1_memCtrl_cacheOpType;
  reg                 entries_1_memCtrl_isPrefetch;
  reg        [31:0]   entries_1_imm;
  reg                 entries_1_usePc;
  reg        [31:0]   entries_1_pcData;
  reg        [3:0]    entries_2_robPtr;
  reg        [5:0]    entries_2_physDest_idx;
  reg                 entries_2_physDestIsFpr;
  reg                 entries_2_writesToPhysReg;
  reg                 entries_2_useSrc1;
  reg        [31:0]   entries_2_src1Data;
  reg        [5:0]    entries_2_src1Tag;
  reg                 entries_2_src1Ready;
  reg                 entries_2_src1IsFpr;
  reg                 entries_2_useSrc2;
  reg        [31:0]   entries_2_src2Data;
  reg        [5:0]    entries_2_src2Tag;
  reg                 entries_2_src2Ready;
  reg                 entries_2_src2IsFpr;
  reg        [1:0]    entries_2_memCtrl_size;
  reg                 entries_2_memCtrl_isSignedLoad;
  reg                 entries_2_memCtrl_isStore;
  reg                 entries_2_memCtrl_isLoadLinked;
  reg                 entries_2_memCtrl_isStoreCond;
  reg        [4:0]    entries_2_memCtrl_atomicOp;
  reg                 entries_2_memCtrl_isFence;
  reg        [7:0]    entries_2_memCtrl_fenceMode;
  reg                 entries_2_memCtrl_isCacheOp;
  reg        [4:0]    entries_2_memCtrl_cacheOpType;
  reg                 entries_2_memCtrl_isPrefetch;
  reg        [31:0]   entries_2_imm;
  reg                 entries_2_usePc;
  reg        [31:0]   entries_2_pcData;
  reg        [3:0]    entries_3_robPtr;
  reg        [5:0]    entries_3_physDest_idx;
  reg                 entries_3_physDestIsFpr;
  reg                 entries_3_writesToPhysReg;
  reg                 entries_3_useSrc1;
  reg        [31:0]   entries_3_src1Data;
  reg        [5:0]    entries_3_src1Tag;
  reg                 entries_3_src1Ready;
  reg                 entries_3_src1IsFpr;
  reg                 entries_3_useSrc2;
  reg        [31:0]   entries_3_src2Data;
  reg        [5:0]    entries_3_src2Tag;
  reg                 entries_3_src2Ready;
  reg                 entries_3_src2IsFpr;
  reg        [1:0]    entries_3_memCtrl_size;
  reg                 entries_3_memCtrl_isSignedLoad;
  reg                 entries_3_memCtrl_isStore;
  reg                 entries_3_memCtrl_isLoadLinked;
  reg                 entries_3_memCtrl_isStoreCond;
  reg        [4:0]    entries_3_memCtrl_atomicOp;
  reg                 entries_3_memCtrl_isFence;
  reg        [7:0]    entries_3_memCtrl_fenceMode;
  reg                 entries_3_memCtrl_isCacheOp;
  reg        [4:0]    entries_3_memCtrl_cacheOpType;
  reg                 entries_3_memCtrl_isPrefetch;
  reg        [31:0]   entries_3_imm;
  reg                 entries_3_usePc;
  reg        [31:0]   entries_3_pcData;
  reg                 entryValids_0;
  reg                 entryValids_1;
  reg                 entryValids_2;
  reg                 entryValids_3;
  wire                io_issueOut_fire;
  wire                localWakeupValid;
  reg        [3:0]    wokeUpSrc1Mask;
  reg        [3:0]    wokeUpSrc2Mask;
  wire                _zz_when_IssueQueueComponent_l103;
  wire                _zz_when_IssueQueueComponent_l106;
  wire                when_IssueQueueComponent_l103;
  wire                when_IssueQueueComponent_l106;
  wire                when_IssueQueueComponent_l113;
  wire                when_IssueQueueComponent_l116;
  wire                when_IssueQueueComponent_l113_1;
  wire                when_IssueQueueComponent_l116_1;
  wire                when_IssueQueueComponent_l113_2;
  wire                when_IssueQueueComponent_l116_2;
  wire                when_IssueQueueComponent_l113_3;
  wire                when_IssueQueueComponent_l116_3;
  wire                when_IssueQueueComponent_l113_4;
  wire                when_IssueQueueComponent_l116_4;
  wire                _zz_when_IssueQueueComponent_l103_1;
  wire                _zz_when_IssueQueueComponent_l106_1;
  wire                when_IssueQueueComponent_l103_1;
  wire                when_IssueQueueComponent_l106_1;
  wire                when_IssueQueueComponent_l113_5;
  wire                when_IssueQueueComponent_l116_5;
  wire                when_IssueQueueComponent_l113_6;
  wire                when_IssueQueueComponent_l116_6;
  wire                when_IssueQueueComponent_l113_7;
  wire                when_IssueQueueComponent_l116_7;
  wire                when_IssueQueueComponent_l113_8;
  wire                when_IssueQueueComponent_l116_8;
  wire                when_IssueQueueComponent_l113_9;
  wire                when_IssueQueueComponent_l116_9;
  wire                _zz_when_IssueQueueComponent_l103_2;
  wire                _zz_when_IssueQueueComponent_l106_2;
  wire                when_IssueQueueComponent_l103_2;
  wire                when_IssueQueueComponent_l106_2;
  wire                when_IssueQueueComponent_l113_10;
  wire                when_IssueQueueComponent_l116_10;
  wire                when_IssueQueueComponent_l113_11;
  wire                when_IssueQueueComponent_l116_11;
  wire                when_IssueQueueComponent_l113_12;
  wire                when_IssueQueueComponent_l116_12;
  wire                when_IssueQueueComponent_l113_13;
  wire                when_IssueQueueComponent_l116_13;
  wire                when_IssueQueueComponent_l113_14;
  wire                when_IssueQueueComponent_l116_14;
  wire                _zz_when_IssueQueueComponent_l103_3;
  wire                _zz_when_IssueQueueComponent_l106_3;
  wire                when_IssueQueueComponent_l103_3;
  wire                when_IssueQueueComponent_l106_3;
  wire                when_IssueQueueComponent_l113_15;
  wire                when_IssueQueueComponent_l116_15;
  wire                when_IssueQueueComponent_l113_16;
  wire                when_IssueQueueComponent_l116_16;
  wire                when_IssueQueueComponent_l113_17;
  wire                when_IssueQueueComponent_l116_17;
  wire                when_IssueQueueComponent_l113_18;
  wire                when_IssueQueueComponent_l116_18;
  wire                when_IssueQueueComponent_l113_19;
  wire                when_IssueQueueComponent_l116_19;
  wire                entriesReadyToIssue_0;
  wire                entriesReadyToIssue_1;
  wire                entriesReadyToIssue_2;
  wire                entriesReadyToIssue_3;
  wire       [3:0]    issueRequestMask;
  wire       [3:0]    issueRequestMask_ohFirst_input;
  wire       [3:0]    issueRequestMask_ohFirst_masked;
  wire       [3:0]    issueRequestOh;
  wire                _zz_issueIdx;
  wire                _zz_issueIdx_1;
  wire                _zz_issueIdx_2;
  wire       [1:0]    issueIdx;
  wire       [1:0]    _zz_io_issueOut_payload_memCtrl_size;
  wire       [3:0]    freeSlotsMask;
  wire                hasSpaceForNewEntry;
  reg        [3:0]    firedSlotMask;
  wire       [3:0]    _zz_allocationMask;
  wire       [3:0]    allocationMask;
  wire                _zz_allocateIdx;
  wire                _zz_allocateIdx_1;
  wire                _zz_allocateIdx_2;
  wire       [1:0]    allocateIdx;
  reg        [3:0]    entriesNext_0_robPtr;
  reg        [5:0]    entriesNext_0_physDest_idx;
  reg                 entriesNext_0_physDestIsFpr;
  reg                 entriesNext_0_writesToPhysReg;
  reg                 entriesNext_0_useSrc1;
  reg        [31:0]   entriesNext_0_src1Data;
  reg        [5:0]    entriesNext_0_src1Tag;
  reg                 entriesNext_0_src1Ready;
  reg                 entriesNext_0_src1IsFpr;
  reg                 entriesNext_0_useSrc2;
  reg        [31:0]   entriesNext_0_src2Data;
  reg        [5:0]    entriesNext_0_src2Tag;
  reg                 entriesNext_0_src2Ready;
  reg                 entriesNext_0_src2IsFpr;
  reg        [1:0]    entriesNext_0_memCtrl_size;
  reg                 entriesNext_0_memCtrl_isSignedLoad;
  reg                 entriesNext_0_memCtrl_isStore;
  reg                 entriesNext_0_memCtrl_isLoadLinked;
  reg                 entriesNext_0_memCtrl_isStoreCond;
  reg        [4:0]    entriesNext_0_memCtrl_atomicOp;
  reg                 entriesNext_0_memCtrl_isFence;
  reg        [7:0]    entriesNext_0_memCtrl_fenceMode;
  reg                 entriesNext_0_memCtrl_isCacheOp;
  reg        [4:0]    entriesNext_0_memCtrl_cacheOpType;
  reg                 entriesNext_0_memCtrl_isPrefetch;
  reg        [31:0]   entriesNext_0_imm;
  reg                 entriesNext_0_usePc;
  reg        [31:0]   entriesNext_0_pcData;
  reg        [3:0]    entriesNext_1_robPtr;
  reg        [5:0]    entriesNext_1_physDest_idx;
  reg                 entriesNext_1_physDestIsFpr;
  reg                 entriesNext_1_writesToPhysReg;
  reg                 entriesNext_1_useSrc1;
  reg        [31:0]   entriesNext_1_src1Data;
  reg        [5:0]    entriesNext_1_src1Tag;
  reg                 entriesNext_1_src1Ready;
  reg                 entriesNext_1_src1IsFpr;
  reg                 entriesNext_1_useSrc2;
  reg        [31:0]   entriesNext_1_src2Data;
  reg        [5:0]    entriesNext_1_src2Tag;
  reg                 entriesNext_1_src2Ready;
  reg                 entriesNext_1_src2IsFpr;
  reg        [1:0]    entriesNext_1_memCtrl_size;
  reg                 entriesNext_1_memCtrl_isSignedLoad;
  reg                 entriesNext_1_memCtrl_isStore;
  reg                 entriesNext_1_memCtrl_isLoadLinked;
  reg                 entriesNext_1_memCtrl_isStoreCond;
  reg        [4:0]    entriesNext_1_memCtrl_atomicOp;
  reg                 entriesNext_1_memCtrl_isFence;
  reg        [7:0]    entriesNext_1_memCtrl_fenceMode;
  reg                 entriesNext_1_memCtrl_isCacheOp;
  reg        [4:0]    entriesNext_1_memCtrl_cacheOpType;
  reg                 entriesNext_1_memCtrl_isPrefetch;
  reg        [31:0]   entriesNext_1_imm;
  reg                 entriesNext_1_usePc;
  reg        [31:0]   entriesNext_1_pcData;
  reg        [3:0]    entriesNext_2_robPtr;
  reg        [5:0]    entriesNext_2_physDest_idx;
  reg                 entriesNext_2_physDestIsFpr;
  reg                 entriesNext_2_writesToPhysReg;
  reg                 entriesNext_2_useSrc1;
  reg        [31:0]   entriesNext_2_src1Data;
  reg        [5:0]    entriesNext_2_src1Tag;
  reg                 entriesNext_2_src1Ready;
  reg                 entriesNext_2_src1IsFpr;
  reg                 entriesNext_2_useSrc2;
  reg        [31:0]   entriesNext_2_src2Data;
  reg        [5:0]    entriesNext_2_src2Tag;
  reg                 entriesNext_2_src2Ready;
  reg                 entriesNext_2_src2IsFpr;
  reg        [1:0]    entriesNext_2_memCtrl_size;
  reg                 entriesNext_2_memCtrl_isSignedLoad;
  reg                 entriesNext_2_memCtrl_isStore;
  reg                 entriesNext_2_memCtrl_isLoadLinked;
  reg                 entriesNext_2_memCtrl_isStoreCond;
  reg        [4:0]    entriesNext_2_memCtrl_atomicOp;
  reg                 entriesNext_2_memCtrl_isFence;
  reg        [7:0]    entriesNext_2_memCtrl_fenceMode;
  reg                 entriesNext_2_memCtrl_isCacheOp;
  reg        [4:0]    entriesNext_2_memCtrl_cacheOpType;
  reg                 entriesNext_2_memCtrl_isPrefetch;
  reg        [31:0]   entriesNext_2_imm;
  reg                 entriesNext_2_usePc;
  reg        [31:0]   entriesNext_2_pcData;
  reg        [3:0]    entriesNext_3_robPtr;
  reg        [5:0]    entriesNext_3_physDest_idx;
  reg                 entriesNext_3_physDestIsFpr;
  reg                 entriesNext_3_writesToPhysReg;
  reg                 entriesNext_3_useSrc1;
  reg        [31:0]   entriesNext_3_src1Data;
  reg        [5:0]    entriesNext_3_src1Tag;
  reg                 entriesNext_3_src1Ready;
  reg                 entriesNext_3_src1IsFpr;
  reg                 entriesNext_3_useSrc2;
  reg        [31:0]   entriesNext_3_src2Data;
  reg        [5:0]    entriesNext_3_src2Tag;
  reg                 entriesNext_3_src2Ready;
  reg                 entriesNext_3_src2IsFpr;
  reg        [1:0]    entriesNext_3_memCtrl_size;
  reg                 entriesNext_3_memCtrl_isSignedLoad;
  reg                 entriesNext_3_memCtrl_isStore;
  reg                 entriesNext_3_memCtrl_isLoadLinked;
  reg                 entriesNext_3_memCtrl_isStoreCond;
  reg        [4:0]    entriesNext_3_memCtrl_atomicOp;
  reg                 entriesNext_3_memCtrl_isFence;
  reg        [7:0]    entriesNext_3_memCtrl_fenceMode;
  reg                 entriesNext_3_memCtrl_isCacheOp;
  reg        [4:0]    entriesNext_3_memCtrl_cacheOpType;
  reg                 entriesNext_3_memCtrl_isPrefetch;
  reg        [31:0]   entriesNext_3_imm;
  reg                 entriesNext_3_usePc;
  reg        [31:0]   entriesNext_3_pcData;
  reg                 entryValidsNext_0;
  reg                 entryValidsNext_1;
  reg                 entryValidsNext_2;
  reg                 entryValidsNext_3;
  wire                when_IssueQueueComponent_l186;
  wire                when_IssueQueueComponent_l187;
  wire                when_IssueQueueComponent_l186_1;
  wire                when_IssueQueueComponent_l187_1;
  wire                when_IssueQueueComponent_l186_2;
  wire                when_IssueQueueComponent_l187_2;
  wire                when_IssueQueueComponent_l186_3;
  wire                when_IssueQueueComponent_l187_3;
  wire       [3:0]    _zz_1;
  wire                io_allocateIn_fire;
  wire       [3:0]    _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_entriesNext_0_src1Ready;
  wire                _zz_entriesNext_0_src2Ready;
  wire       [3:0]    _zz_7;
  wire                when_IssueQueueComponent_l212;
  wire                when_IssueQueueComponent_l215;
  wire                when_IssueQueueComponent_l212_1;
  wire                when_IssueQueueComponent_l215_1;
  wire                when_IssueQueueComponent_l212_2;
  wire                when_IssueQueueComponent_l215_2;
  wire                when_IssueQueueComponent_l212_3;
  wire                when_IssueQueueComponent_l215_3;
  wire                when_IssueQueueComponent_l212_4;
  wire                when_IssueQueueComponent_l215_4;
  wire       [2:0]    _zz_currentValidCount;
  wire       [2:0]    _zz_currentValidCount_1;
  wire       [2:0]    _zz_currentValidCount_2;
  wire       [2:0]    _zz_currentValidCount_3;
  wire       [2:0]    _zz_currentValidCount_4;
  wire       [2:0]    _zz_currentValidCount_5;
  wire       [2:0]    _zz_currentValidCount_6;
  wire       [2:0]    _zz_currentValidCount_7;
  wire       [2:0]    currentValidCount;
  wire                logCondition;
  wire                when_IssueQueueComponent_l256;
  `ifndef SYNTHESIS
  reg [87:0] io_allocateIn_payload_uop_decoded_uopCode_string;
  reg [151:0] io_allocateIn_payload_uop_decoded_exeUnit_string;
  reg [71:0] io_allocateIn_payload_uop_decoded_isa_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] io_allocateIn_payload_uop_decoded_immUsage_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] io_allocateIn_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_allocateIn_payload_uop_decoded_decodeExceptionCode_string;
  reg [7:0] io_issueOut_payload_memCtrl_size_string;
  reg [7:0] entries_0_memCtrl_size_string;
  reg [7:0] entries_1_memCtrl_size_string;
  reg [7:0] entries_2_memCtrl_size_string;
  reg [7:0] entries_3_memCtrl_size_string;
  reg [7:0] _zz_io_issueOut_payload_memCtrl_size_string;
  reg [7:0] entriesNext_0_memCtrl_size_string;
  reg [7:0] entriesNext_1_memCtrl_size_string;
  reg [7:0] entriesNext_2_memCtrl_size_string;
  reg [7:0] entriesNext_3_memCtrl_size_string;
  `endif


  assign _zz_issueRequestMask_ohFirst_masked = (issueRequestMask_ohFirst_input - 4'b0001);
  assign _zz_allocationMask_1 = (_zz_allocationMask - 4'b0001);
  assign _zz_currentValidCount_12 = entryValids_3;
  assign _zz_currentValidCount_11 = {2'd0, _zz_currentValidCount_12};
  assign _zz_currentValidCount_9 = {entryValids_2,{entryValids_1,entryValids_0}};
  always @(*) begin
    case(issueIdx)
      2'b00 : begin
        _zz__zz_io_issueOut_payload_memCtrl_size = entries_0_memCtrl_size;
        _zz_io_issueOut_payload_robPtr = entries_0_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_0_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_0_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_0_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_0_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_0_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_0_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_0_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_0_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_0_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_0_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_0_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_0_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_0_src2IsFpr;
        _zz_io_issueOut_payload_memCtrl_isSignedLoad = entries_0_memCtrl_isSignedLoad;
        _zz_io_issueOut_payload_memCtrl_isStore = entries_0_memCtrl_isStore;
        _zz_io_issueOut_payload_memCtrl_isLoadLinked = entries_0_memCtrl_isLoadLinked;
        _zz_io_issueOut_payload_memCtrl_isStoreCond = entries_0_memCtrl_isStoreCond;
        _zz_io_issueOut_payload_memCtrl_atomicOp = entries_0_memCtrl_atomicOp;
        _zz_io_issueOut_payload_memCtrl_isFence = entries_0_memCtrl_isFence;
        _zz_io_issueOut_payload_memCtrl_fenceMode = entries_0_memCtrl_fenceMode;
        _zz_io_issueOut_payload_memCtrl_isCacheOp = entries_0_memCtrl_isCacheOp;
        _zz_io_issueOut_payload_memCtrl_cacheOpType = entries_0_memCtrl_cacheOpType;
        _zz_io_issueOut_payload_memCtrl_isPrefetch = entries_0_memCtrl_isPrefetch;
        _zz_io_issueOut_payload_imm = entries_0_imm;
        _zz_io_issueOut_payload_usePc = entries_0_usePc;
        _zz_io_issueOut_payload_pcData = entries_0_pcData;
      end
      2'b01 : begin
        _zz__zz_io_issueOut_payload_memCtrl_size = entries_1_memCtrl_size;
        _zz_io_issueOut_payload_robPtr = entries_1_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_1_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_1_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_1_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_1_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_1_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_1_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_1_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_1_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_1_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_1_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_1_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_1_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_1_src2IsFpr;
        _zz_io_issueOut_payload_memCtrl_isSignedLoad = entries_1_memCtrl_isSignedLoad;
        _zz_io_issueOut_payload_memCtrl_isStore = entries_1_memCtrl_isStore;
        _zz_io_issueOut_payload_memCtrl_isLoadLinked = entries_1_memCtrl_isLoadLinked;
        _zz_io_issueOut_payload_memCtrl_isStoreCond = entries_1_memCtrl_isStoreCond;
        _zz_io_issueOut_payload_memCtrl_atomicOp = entries_1_memCtrl_atomicOp;
        _zz_io_issueOut_payload_memCtrl_isFence = entries_1_memCtrl_isFence;
        _zz_io_issueOut_payload_memCtrl_fenceMode = entries_1_memCtrl_fenceMode;
        _zz_io_issueOut_payload_memCtrl_isCacheOp = entries_1_memCtrl_isCacheOp;
        _zz_io_issueOut_payload_memCtrl_cacheOpType = entries_1_memCtrl_cacheOpType;
        _zz_io_issueOut_payload_memCtrl_isPrefetch = entries_1_memCtrl_isPrefetch;
        _zz_io_issueOut_payload_imm = entries_1_imm;
        _zz_io_issueOut_payload_usePc = entries_1_usePc;
        _zz_io_issueOut_payload_pcData = entries_1_pcData;
      end
      2'b10 : begin
        _zz__zz_io_issueOut_payload_memCtrl_size = entries_2_memCtrl_size;
        _zz_io_issueOut_payload_robPtr = entries_2_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_2_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_2_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_2_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_2_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_2_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_2_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_2_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_2_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_2_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_2_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_2_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_2_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_2_src2IsFpr;
        _zz_io_issueOut_payload_memCtrl_isSignedLoad = entries_2_memCtrl_isSignedLoad;
        _zz_io_issueOut_payload_memCtrl_isStore = entries_2_memCtrl_isStore;
        _zz_io_issueOut_payload_memCtrl_isLoadLinked = entries_2_memCtrl_isLoadLinked;
        _zz_io_issueOut_payload_memCtrl_isStoreCond = entries_2_memCtrl_isStoreCond;
        _zz_io_issueOut_payload_memCtrl_atomicOp = entries_2_memCtrl_atomicOp;
        _zz_io_issueOut_payload_memCtrl_isFence = entries_2_memCtrl_isFence;
        _zz_io_issueOut_payload_memCtrl_fenceMode = entries_2_memCtrl_fenceMode;
        _zz_io_issueOut_payload_memCtrl_isCacheOp = entries_2_memCtrl_isCacheOp;
        _zz_io_issueOut_payload_memCtrl_cacheOpType = entries_2_memCtrl_cacheOpType;
        _zz_io_issueOut_payload_memCtrl_isPrefetch = entries_2_memCtrl_isPrefetch;
        _zz_io_issueOut_payload_imm = entries_2_imm;
        _zz_io_issueOut_payload_usePc = entries_2_usePc;
        _zz_io_issueOut_payload_pcData = entries_2_pcData;
      end
      default : begin
        _zz__zz_io_issueOut_payload_memCtrl_size = entries_3_memCtrl_size;
        _zz_io_issueOut_payload_robPtr = entries_3_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_3_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_3_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_3_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_3_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_3_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_3_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_3_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_3_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_3_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_3_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_3_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_3_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_3_src2IsFpr;
        _zz_io_issueOut_payload_memCtrl_isSignedLoad = entries_3_memCtrl_isSignedLoad;
        _zz_io_issueOut_payload_memCtrl_isStore = entries_3_memCtrl_isStore;
        _zz_io_issueOut_payload_memCtrl_isLoadLinked = entries_3_memCtrl_isLoadLinked;
        _zz_io_issueOut_payload_memCtrl_isStoreCond = entries_3_memCtrl_isStoreCond;
        _zz_io_issueOut_payload_memCtrl_atomicOp = entries_3_memCtrl_atomicOp;
        _zz_io_issueOut_payload_memCtrl_isFence = entries_3_memCtrl_isFence;
        _zz_io_issueOut_payload_memCtrl_fenceMode = entries_3_memCtrl_fenceMode;
        _zz_io_issueOut_payload_memCtrl_isCacheOp = entries_3_memCtrl_isCacheOp;
        _zz_io_issueOut_payload_memCtrl_cacheOpType = entries_3_memCtrl_cacheOpType;
        _zz_io_issueOut_payload_memCtrl_isPrefetch = entries_3_memCtrl_isPrefetch;
        _zz_io_issueOut_payload_imm = entries_3_imm;
        _zz_io_issueOut_payload_usePc = entries_3_usePc;
        _zz_io_issueOut_payload_pcData = entries_3_pcData;
      end
    endcase
  end

  always @(*) begin
    case(_zz_currentValidCount_9)
      3'b000 : _zz_currentValidCount_8 = _zz_currentValidCount;
      3'b001 : _zz_currentValidCount_8 = _zz_currentValidCount_1;
      3'b010 : _zz_currentValidCount_8 = _zz_currentValidCount_2;
      3'b011 : _zz_currentValidCount_8 = _zz_currentValidCount_3;
      3'b100 : _zz_currentValidCount_8 = _zz_currentValidCount_4;
      3'b101 : _zz_currentValidCount_8 = _zz_currentValidCount_5;
      3'b110 : _zz_currentValidCount_8 = _zz_currentValidCount_6;
      default : _zz_currentValidCount_8 = _zz_currentValidCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_currentValidCount_11)
      3'b000 : _zz_currentValidCount_10 = _zz_currentValidCount;
      3'b001 : _zz_currentValidCount_10 = _zz_currentValidCount_1;
      3'b010 : _zz_currentValidCount_10 = _zz_currentValidCount_2;
      3'b011 : _zz_currentValidCount_10 = _zz_currentValidCount_3;
      3'b100 : _zz_currentValidCount_10 = _zz_currentValidCount_4;
      3'b101 : _zz_currentValidCount_10 = _zz_currentValidCount_5;
      3'b110 : _zz_currentValidCount_10 = _zz_currentValidCount_6;
      default : _zz_currentValidCount_10 = _zz_currentValidCount_7;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : io_allocateIn_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_allocateIn_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_allocateIn_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_allocateIn_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_allocateIn_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_allocateIn_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_allocateIn_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_allocateIn_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_allocateIn_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_allocateIn_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_allocateIn_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_allocateIn_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_allocateIn_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_allocateIn_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_allocateIn_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_allocateIn_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_allocateIn_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : io_allocateIn_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : io_allocateIn_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_allocateIn_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_allocateIn_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_allocateIn_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_allocateIn_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_allocateIn_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_allocateIn_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_isa)
      IsaType_UNKNOWN : io_allocateIn_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_allocateIn_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : io_allocateIn_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_allocateIn_payload_uop_decoded_isa_string = "LOONGARCH";
      default : io_allocateIn_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : io_allocateIn_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : io_allocateIn_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "D";
      default : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_memCtrl_size)
      MemAccessSize_B : io_issueOut_payload_memCtrl_size_string = "B";
      MemAccessSize_H : io_issueOut_payload_memCtrl_size_string = "H";
      MemAccessSize_W : io_issueOut_payload_memCtrl_size_string = "W";
      MemAccessSize_D : io_issueOut_payload_memCtrl_size_string = "D";
      default : io_issueOut_payload_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_0_memCtrl_size)
      MemAccessSize_B : entries_0_memCtrl_size_string = "B";
      MemAccessSize_H : entries_0_memCtrl_size_string = "H";
      MemAccessSize_W : entries_0_memCtrl_size_string = "W";
      MemAccessSize_D : entries_0_memCtrl_size_string = "D";
      default : entries_0_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_1_memCtrl_size)
      MemAccessSize_B : entries_1_memCtrl_size_string = "B";
      MemAccessSize_H : entries_1_memCtrl_size_string = "H";
      MemAccessSize_W : entries_1_memCtrl_size_string = "W";
      MemAccessSize_D : entries_1_memCtrl_size_string = "D";
      default : entries_1_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_2_memCtrl_size)
      MemAccessSize_B : entries_2_memCtrl_size_string = "B";
      MemAccessSize_H : entries_2_memCtrl_size_string = "H";
      MemAccessSize_W : entries_2_memCtrl_size_string = "W";
      MemAccessSize_D : entries_2_memCtrl_size_string = "D";
      default : entries_2_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_3_memCtrl_size)
      MemAccessSize_B : entries_3_memCtrl_size_string = "B";
      MemAccessSize_H : entries_3_memCtrl_size_string = "H";
      MemAccessSize_W : entries_3_memCtrl_size_string = "W";
      MemAccessSize_D : entries_3_memCtrl_size_string = "D";
      default : entries_3_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_memCtrl_size)
      MemAccessSize_B : _zz_io_issueOut_payload_memCtrl_size_string = "B";
      MemAccessSize_H : _zz_io_issueOut_payload_memCtrl_size_string = "H";
      MemAccessSize_W : _zz_io_issueOut_payload_memCtrl_size_string = "W";
      MemAccessSize_D : _zz_io_issueOut_payload_memCtrl_size_string = "D";
      default : _zz_io_issueOut_payload_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_memCtrl_size)
      MemAccessSize_B : entriesNext_0_memCtrl_size_string = "B";
      MemAccessSize_H : entriesNext_0_memCtrl_size_string = "H";
      MemAccessSize_W : entriesNext_0_memCtrl_size_string = "W";
      MemAccessSize_D : entriesNext_0_memCtrl_size_string = "D";
      default : entriesNext_0_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_memCtrl_size)
      MemAccessSize_B : entriesNext_1_memCtrl_size_string = "B";
      MemAccessSize_H : entriesNext_1_memCtrl_size_string = "H";
      MemAccessSize_W : entriesNext_1_memCtrl_size_string = "W";
      MemAccessSize_D : entriesNext_1_memCtrl_size_string = "D";
      default : entriesNext_1_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_memCtrl_size)
      MemAccessSize_B : entriesNext_2_memCtrl_size_string = "B";
      MemAccessSize_H : entriesNext_2_memCtrl_size_string = "H";
      MemAccessSize_W : entriesNext_2_memCtrl_size_string = "W";
      MemAccessSize_D : entriesNext_2_memCtrl_size_string = "D";
      default : entriesNext_2_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_memCtrl_size)
      MemAccessSize_B : entriesNext_3_memCtrl_size_string = "B";
      MemAccessSize_H : entriesNext_3_memCtrl_size_string = "H";
      MemAccessSize_W : entriesNext_3_memCtrl_size_string = "W";
      MemAccessSize_D : entriesNext_3_memCtrl_size_string = "D";
      default : entriesNext_3_memCtrl_size_string = "?";
    endcase
  end
  `endif

  assign io_issueOut_fire = (io_issueOut_valid && io_issueOut_ready);
  assign localWakeupValid = (io_issueOut_fire && io_issueOut_payload_writesToPhysReg);
  always @(*) begin
    wokeUpSrc1Mask = 4'b0000;
    if(entryValids_0) begin
      if(when_IssueQueueComponent_l103) begin
        wokeUpSrc1Mask[0] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_1) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_2) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_3) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_4) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
    end
    if(entryValids_1) begin
      if(when_IssueQueueComponent_l103_1) begin
        wokeUpSrc1Mask[1] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_5) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_6) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_7) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_8) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_9) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
    end
    if(entryValids_2) begin
      if(when_IssueQueueComponent_l103_2) begin
        wokeUpSrc1Mask[2] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_10) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_11) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_12) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_13) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_14) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
    end
    if(entryValids_3) begin
      if(when_IssueQueueComponent_l103_3) begin
        wokeUpSrc1Mask[3] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_15) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_16) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_17) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_18) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_19) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    wokeUpSrc2Mask = 4'b0000;
    if(entryValids_0) begin
      if(when_IssueQueueComponent_l106) begin
        wokeUpSrc2Mask[0] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_1) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_2) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_3) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_4) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
    end
    if(entryValids_1) begin
      if(when_IssueQueueComponent_l106_1) begin
        wokeUpSrc2Mask[1] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_5) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_6) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_7) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_8) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_9) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
    end
    if(entryValids_2) begin
      if(when_IssueQueueComponent_l106_2) begin
        wokeUpSrc2Mask[2] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_10) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_11) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_12) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_13) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_14) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
    end
    if(entryValids_3) begin
      if(when_IssueQueueComponent_l106_3) begin
        wokeUpSrc2Mask[3] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_15) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_16) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_17) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_18) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_19) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
    end
  end

  assign _zz_when_IssueQueueComponent_l103 = ((! entries_0_src1Ready) && entries_0_useSrc1);
  assign _zz_when_IssueQueueComponent_l106 = ((! entries_0_src2Ready) && entries_0_useSrc2);
  assign when_IssueQueueComponent_l103 = ((_zz_when_IssueQueueComponent_l103 && localWakeupValid) && (entries_0_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106 = ((_zz_when_IssueQueueComponent_l106 && localWakeupValid) && (entries_0_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_1 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_1 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_2 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_2 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_3 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_3 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_4 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_4 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_1 = ((! entries_1_src1Ready) && entries_1_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_1 = ((! entries_1_src2Ready) && entries_1_useSrc2);
  assign when_IssueQueueComponent_l103_1 = ((_zz_when_IssueQueueComponent_l103_1 && localWakeupValid) && (entries_1_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_1 = ((_zz_when_IssueQueueComponent_l106_1 && localWakeupValid) && (entries_1_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_5 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_5 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_6 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_6 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_7 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_7 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_8 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_8 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_9 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_9 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_2 = ((! entries_2_src1Ready) && entries_2_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_2 = ((! entries_2_src2Ready) && entries_2_useSrc2);
  assign when_IssueQueueComponent_l103_2 = ((_zz_when_IssueQueueComponent_l103_2 && localWakeupValid) && (entries_2_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_2 = ((_zz_when_IssueQueueComponent_l106_2 && localWakeupValid) && (entries_2_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_10 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_10 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_11 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_11 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_12 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_12 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_13 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_13 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_14 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_14 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_3 = ((! entries_3_src1Ready) && entries_3_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_3 = ((! entries_3_src2Ready) && entries_3_useSrc2);
  assign when_IssueQueueComponent_l103_3 = ((_zz_when_IssueQueueComponent_l103_3 && localWakeupValid) && (entries_3_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_3 = ((_zz_when_IssueQueueComponent_l106_3 && localWakeupValid) && (entries_3_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_15 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_15 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_16 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_16 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_17 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_17 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_18 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_18 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_19 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_19 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign entriesReadyToIssue_0 = ((entryValids_0 && ((! entries_0_useSrc1) || entries_0_src1Ready)) && ((! entries_0_useSrc2) || entries_0_src2Ready));
  assign entriesReadyToIssue_1 = ((entryValids_1 && ((! entries_1_useSrc1) || entries_1_src1Ready)) && ((! entries_1_useSrc2) || entries_1_src2Ready));
  assign entriesReadyToIssue_2 = ((entryValids_2 && ((! entries_2_useSrc1) || entries_2_src1Ready)) && ((! entries_2_useSrc2) || entries_2_src2Ready));
  assign entriesReadyToIssue_3 = ((entryValids_3 && ((! entries_3_useSrc1) || entries_3_src1Ready)) && ((! entries_3_useSrc2) || entries_3_src2Ready));
  assign issueRequestMask = {entriesReadyToIssue_3,{entriesReadyToIssue_2,{entriesReadyToIssue_1,entriesReadyToIssue_0}}};
  assign issueRequestMask_ohFirst_input = issueRequestMask;
  assign issueRequestMask_ohFirst_masked = (issueRequestMask_ohFirst_input & (~ _zz_issueRequestMask_ohFirst_masked));
  assign issueRequestOh = issueRequestMask_ohFirst_masked;
  assign _zz_issueIdx = issueRequestOh[3];
  assign _zz_issueIdx_1 = (issueRequestOh[1] || _zz_issueIdx);
  assign _zz_issueIdx_2 = (issueRequestOh[2] || _zz_issueIdx);
  assign issueIdx = {_zz_issueIdx_2,_zz_issueIdx_1};
  assign io_issueOut_valid = ((|issueRequestOh) && (! io_flush));
  assign _zz_io_issueOut_payload_memCtrl_size = _zz__zz_io_issueOut_payload_memCtrl_size;
  assign io_issueOut_payload_robPtr = _zz_io_issueOut_payload_robPtr;
  assign io_issueOut_payload_physDest_idx = _zz_io_issueOut_payload_physDest_idx;
  assign io_issueOut_payload_physDestIsFpr = _zz_io_issueOut_payload_physDestIsFpr;
  assign io_issueOut_payload_writesToPhysReg = _zz_io_issueOut_payload_writesToPhysReg;
  assign io_issueOut_payload_useSrc1 = _zz_io_issueOut_payload_useSrc1;
  assign io_issueOut_payload_src1Data = _zz_io_issueOut_payload_src1Data;
  assign io_issueOut_payload_src1Tag = _zz_io_issueOut_payload_src1Tag;
  assign io_issueOut_payload_src1Ready = _zz_io_issueOut_payload_src1Ready;
  assign io_issueOut_payload_src1IsFpr = _zz_io_issueOut_payload_src1IsFpr;
  assign io_issueOut_payload_useSrc2 = _zz_io_issueOut_payload_useSrc2;
  assign io_issueOut_payload_src2Data = _zz_io_issueOut_payload_src2Data;
  assign io_issueOut_payload_src2Tag = _zz_io_issueOut_payload_src2Tag;
  assign io_issueOut_payload_src2Ready = _zz_io_issueOut_payload_src2Ready;
  assign io_issueOut_payload_src2IsFpr = _zz_io_issueOut_payload_src2IsFpr;
  assign io_issueOut_payload_memCtrl_size = _zz_io_issueOut_payload_memCtrl_size;
  assign io_issueOut_payload_memCtrl_isSignedLoad = _zz_io_issueOut_payload_memCtrl_isSignedLoad;
  assign io_issueOut_payload_memCtrl_isStore = _zz_io_issueOut_payload_memCtrl_isStore;
  assign io_issueOut_payload_memCtrl_isLoadLinked = _zz_io_issueOut_payload_memCtrl_isLoadLinked;
  assign io_issueOut_payload_memCtrl_isStoreCond = _zz_io_issueOut_payload_memCtrl_isStoreCond;
  assign io_issueOut_payload_memCtrl_atomicOp = _zz_io_issueOut_payload_memCtrl_atomicOp;
  assign io_issueOut_payload_memCtrl_isFence = _zz_io_issueOut_payload_memCtrl_isFence;
  assign io_issueOut_payload_memCtrl_fenceMode = _zz_io_issueOut_payload_memCtrl_fenceMode;
  assign io_issueOut_payload_memCtrl_isCacheOp = _zz_io_issueOut_payload_memCtrl_isCacheOp;
  assign io_issueOut_payload_memCtrl_cacheOpType = _zz_io_issueOut_payload_memCtrl_cacheOpType;
  assign io_issueOut_payload_memCtrl_isPrefetch = _zz_io_issueOut_payload_memCtrl_isPrefetch;
  assign io_issueOut_payload_imm = _zz_io_issueOut_payload_imm;
  assign io_issueOut_payload_usePc = _zz_io_issueOut_payload_usePc;
  assign io_issueOut_payload_pcData = _zz_io_issueOut_payload_pcData;
  assign freeSlotsMask = {(! entryValids_3),{(! entryValids_2),{(! entryValids_1),(! entryValids_0)}}};
  assign hasSpaceForNewEntry = ((|freeSlotsMask) || io_issueOut_fire);
  assign io_allocateIn_ready = (hasSpaceForNewEntry && (! io_flush));
  always @(*) begin
    firedSlotMask = 4'b0000;
    if(io_issueOut_fire) begin
      firedSlotMask[issueIdx] = 1'b1;
    end
  end

  assign _zz_allocationMask = (freeSlotsMask | firedSlotMask);
  assign allocationMask = (_zz_allocationMask & (~ _zz_allocationMask_1));
  assign _zz_allocateIdx = allocationMask[3];
  assign _zz_allocateIdx_1 = (allocationMask[1] || _zz_allocateIdx);
  assign _zz_allocateIdx_2 = (allocationMask[2] || _zz_allocateIdx);
  assign allocateIdx = {_zz_allocateIdx_2,_zz_allocateIdx_1};
  always @(*) begin
    entriesNext_0_robPtr = entries_0_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_physDest_idx = entries_0_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_physDestIsFpr = entries_0_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_writesToPhysReg = entries_0_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_0_useSrc1 = entries_0_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Data = entries_0_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Tag = entries_0_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Ready = entries_0_src1Ready;
    if(when_IssueQueueComponent_l186) begin
      entriesNext_0_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_3) begin
        entriesNext_0_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1IsFpr = entries_0_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_useSrc2 = entries_0_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Data = entries_0_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Tag = entries_0_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Ready = entries_0_src2Ready;
    if(when_IssueQueueComponent_l187) begin
      entriesNext_0_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_3) begin
        entriesNext_0_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2IsFpr = entries_0_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_size = entries_0_memCtrl_size;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_size = io_allocateIn_payload_uop_decoded_memCtrl_size;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_isSignedLoad = entries_0_memCtrl_isSignedLoad;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_isSignedLoad = io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_isStore = entries_0_memCtrl_isStore;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_isStore = io_allocateIn_payload_uop_decoded_memCtrl_isStore;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_isLoadLinked = entries_0_memCtrl_isLoadLinked;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_isLoadLinked = io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_isStoreCond = entries_0_memCtrl_isStoreCond;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_isStoreCond = io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_atomicOp = entries_0_memCtrl_atomicOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_atomicOp = io_allocateIn_payload_uop_decoded_memCtrl_atomicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_isFence = entries_0_memCtrl_isFence;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_isFence = io_allocateIn_payload_uop_decoded_memCtrl_isFence;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_fenceMode = entries_0_memCtrl_fenceMode;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_fenceMode = io_allocateIn_payload_uop_decoded_memCtrl_fenceMode;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_isCacheOp = entries_0_memCtrl_isCacheOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_isCacheOp = io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_cacheOpType = entries_0_memCtrl_cacheOpType;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_cacheOpType = io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_0_memCtrl_isPrefetch = entries_0_memCtrl_isPrefetch;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_memCtrl_isPrefetch = io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch;
      end
    end
  end

  always @(*) begin
    entriesNext_0_imm = entries_0_imm;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_0_usePc = entries_0_usePc;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_usePc = io_allocateIn_payload_uop_decoded_usePcForAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_pcData = entries_0_pcData;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_pcData = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_1_robPtr = entries_1_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_physDest_idx = entries_1_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_physDestIsFpr = entries_1_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_writesToPhysReg = entries_1_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_1_useSrc1 = entries_1_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Data = entries_1_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Tag = entries_1_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Ready = entries_1_src1Ready;
    if(when_IssueQueueComponent_l186_1) begin
      entriesNext_1_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_4) begin
        entriesNext_1_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1IsFpr = entries_1_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_useSrc2 = entries_1_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Data = entries_1_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Tag = entries_1_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Ready = entries_1_src2Ready;
    if(when_IssueQueueComponent_l187_1) begin
      entriesNext_1_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_4) begin
        entriesNext_1_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2IsFpr = entries_1_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_size = entries_1_memCtrl_size;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_size = io_allocateIn_payload_uop_decoded_memCtrl_size;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_isSignedLoad = entries_1_memCtrl_isSignedLoad;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_isSignedLoad = io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_isStore = entries_1_memCtrl_isStore;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_isStore = io_allocateIn_payload_uop_decoded_memCtrl_isStore;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_isLoadLinked = entries_1_memCtrl_isLoadLinked;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_isLoadLinked = io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_isStoreCond = entries_1_memCtrl_isStoreCond;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_isStoreCond = io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_atomicOp = entries_1_memCtrl_atomicOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_atomicOp = io_allocateIn_payload_uop_decoded_memCtrl_atomicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_isFence = entries_1_memCtrl_isFence;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_isFence = io_allocateIn_payload_uop_decoded_memCtrl_isFence;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_fenceMode = entries_1_memCtrl_fenceMode;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_fenceMode = io_allocateIn_payload_uop_decoded_memCtrl_fenceMode;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_isCacheOp = entries_1_memCtrl_isCacheOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_isCacheOp = io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_cacheOpType = entries_1_memCtrl_cacheOpType;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_cacheOpType = io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_1_memCtrl_isPrefetch = entries_1_memCtrl_isPrefetch;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_memCtrl_isPrefetch = io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch;
      end
    end
  end

  always @(*) begin
    entriesNext_1_imm = entries_1_imm;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_1_usePc = entries_1_usePc;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_usePc = io_allocateIn_payload_uop_decoded_usePcForAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_pcData = entries_1_pcData;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_pcData = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_2_robPtr = entries_2_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_physDest_idx = entries_2_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_physDestIsFpr = entries_2_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_writesToPhysReg = entries_2_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_2_useSrc1 = entries_2_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Data = entries_2_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Tag = entries_2_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Ready = entries_2_src1Ready;
    if(when_IssueQueueComponent_l186_2) begin
      entriesNext_2_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_5) begin
        entriesNext_2_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1IsFpr = entries_2_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_useSrc2 = entries_2_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Data = entries_2_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Tag = entries_2_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Ready = entries_2_src2Ready;
    if(when_IssueQueueComponent_l187_2) begin
      entriesNext_2_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_5) begin
        entriesNext_2_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2IsFpr = entries_2_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_size = entries_2_memCtrl_size;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_size = io_allocateIn_payload_uop_decoded_memCtrl_size;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_isSignedLoad = entries_2_memCtrl_isSignedLoad;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_isSignedLoad = io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_isStore = entries_2_memCtrl_isStore;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_isStore = io_allocateIn_payload_uop_decoded_memCtrl_isStore;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_isLoadLinked = entries_2_memCtrl_isLoadLinked;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_isLoadLinked = io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_isStoreCond = entries_2_memCtrl_isStoreCond;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_isStoreCond = io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_atomicOp = entries_2_memCtrl_atomicOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_atomicOp = io_allocateIn_payload_uop_decoded_memCtrl_atomicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_isFence = entries_2_memCtrl_isFence;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_isFence = io_allocateIn_payload_uop_decoded_memCtrl_isFence;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_fenceMode = entries_2_memCtrl_fenceMode;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_fenceMode = io_allocateIn_payload_uop_decoded_memCtrl_fenceMode;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_isCacheOp = entries_2_memCtrl_isCacheOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_isCacheOp = io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_cacheOpType = entries_2_memCtrl_cacheOpType;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_cacheOpType = io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_2_memCtrl_isPrefetch = entries_2_memCtrl_isPrefetch;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_memCtrl_isPrefetch = io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch;
      end
    end
  end

  always @(*) begin
    entriesNext_2_imm = entries_2_imm;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_2_usePc = entries_2_usePc;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_usePc = io_allocateIn_payload_uop_decoded_usePcForAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_pcData = entries_2_pcData;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_pcData = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_3_robPtr = entries_3_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_physDest_idx = entries_3_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_physDestIsFpr = entries_3_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_writesToPhysReg = entries_3_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_3_useSrc1 = entries_3_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Data = entries_3_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Tag = entries_3_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Ready = entries_3_src1Ready;
    if(when_IssueQueueComponent_l186_3) begin
      entriesNext_3_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_6) begin
        entriesNext_3_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1IsFpr = entries_3_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_useSrc2 = entries_3_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Data = entries_3_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Tag = entries_3_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Ready = entries_3_src2Ready;
    if(when_IssueQueueComponent_l187_3) begin
      entriesNext_3_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_6) begin
        entriesNext_3_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2IsFpr = entries_3_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_size = entries_3_memCtrl_size;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_size = io_allocateIn_payload_uop_decoded_memCtrl_size;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_isSignedLoad = entries_3_memCtrl_isSignedLoad;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_isSignedLoad = io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_isStore = entries_3_memCtrl_isStore;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_isStore = io_allocateIn_payload_uop_decoded_memCtrl_isStore;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_isLoadLinked = entries_3_memCtrl_isLoadLinked;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_isLoadLinked = io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_isStoreCond = entries_3_memCtrl_isStoreCond;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_isStoreCond = io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_atomicOp = entries_3_memCtrl_atomicOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_atomicOp = io_allocateIn_payload_uop_decoded_memCtrl_atomicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_isFence = entries_3_memCtrl_isFence;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_isFence = io_allocateIn_payload_uop_decoded_memCtrl_isFence;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_fenceMode = entries_3_memCtrl_fenceMode;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_fenceMode = io_allocateIn_payload_uop_decoded_memCtrl_fenceMode;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_isCacheOp = entries_3_memCtrl_isCacheOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_isCacheOp = io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_cacheOpType = entries_3_memCtrl_cacheOpType;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_cacheOpType = io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_3_memCtrl_isPrefetch = entries_3_memCtrl_isPrefetch;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_memCtrl_isPrefetch = io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch;
      end
    end
  end

  always @(*) begin
    entriesNext_3_imm = entries_3_imm;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_3_usePc = entries_3_usePc;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_usePc = io_allocateIn_payload_uop_decoded_usePcForAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_pcData = entries_3_pcData;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_pcData = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entryValidsNext_0 = entryValids_0;
    if(io_issueOut_fire) begin
      if(_zz_1[0]) begin
        entryValidsNext_0 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[0]) begin
        entryValidsNext_0 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_0 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_1 = entryValids_1;
    if(io_issueOut_fire) begin
      if(_zz_1[1]) begin
        entryValidsNext_1 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[1]) begin
        entryValidsNext_1 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_1 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_2 = entryValids_2;
    if(io_issueOut_fire) begin
      if(_zz_1[2]) begin
        entryValidsNext_2 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[2]) begin
        entryValidsNext_2 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_2 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_3 = entryValids_3;
    if(io_issueOut_fire) begin
      if(_zz_1[3]) begin
        entryValidsNext_3 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[3]) begin
        entryValidsNext_3 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_3 = 1'b0;
    end
  end

  assign when_IssueQueueComponent_l186 = wokeUpSrc1Mask[0];
  assign when_IssueQueueComponent_l187 = wokeUpSrc2Mask[0];
  assign when_IssueQueueComponent_l186_1 = wokeUpSrc1Mask[1];
  assign when_IssueQueueComponent_l187_1 = wokeUpSrc2Mask[1];
  assign when_IssueQueueComponent_l186_2 = wokeUpSrc1Mask[2];
  assign when_IssueQueueComponent_l187_2 = wokeUpSrc2Mask[2];
  assign when_IssueQueueComponent_l186_3 = wokeUpSrc1Mask[3];
  assign when_IssueQueueComponent_l187_3 = wokeUpSrc2Mask[3];
  assign _zz_1 = ({3'd0,1'b1} <<< issueIdx);
  assign io_allocateIn_fire = (io_allocateIn_valid && io_allocateIn_ready);
  assign _zz_2 = ({3'd0,1'b1} <<< allocateIdx);
  assign _zz_3 = _zz_2[0];
  assign _zz_4 = _zz_2[1];
  assign _zz_5 = _zz_2[2];
  assign _zz_6 = _zz_2[3];
  assign _zz_entriesNext_0_src1Ready = (! io_allocateIn_payload_uop_decoded_useArchSrc1);
  assign _zz_entriesNext_0_src2Ready = (! io_allocateIn_payload_uop_decoded_useArchSrc2);
  assign _zz_7 = ({3'd0,1'b1} <<< allocateIdx);
  assign when_IssueQueueComponent_l212 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l215 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_1 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_1 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_2 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_2 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_3 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_3 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_4 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_4 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_currentValidCount = 3'b000;
  assign _zz_currentValidCount_1 = 3'b001;
  assign _zz_currentValidCount_2 = 3'b001;
  assign _zz_currentValidCount_3 = 3'b010;
  assign _zz_currentValidCount_4 = 3'b001;
  assign _zz_currentValidCount_5 = 3'b010;
  assign _zz_currentValidCount_6 = 3'b010;
  assign _zz_currentValidCount_7 = 3'b011;
  assign currentValidCount = (_zz_currentValidCount_8 + _zz_currentValidCount_10);
  assign logCondition = (io_allocateIn_fire || io_issueOut_fire);
  assign when_IssueQueueComponent_l256 = (logCondition && (3'b000 < currentValidCount));
  always @(posedge clk) begin
    if(reset) begin
      entryValids_0 <= 1'b0;
      entryValids_1 <= 1'b0;
      entryValids_2 <= 1'b0;
      entryValids_3 <= 1'b0;
    end else begin
      entryValids_0 <= entryValidsNext_0;
      entryValids_1 <= entryValidsNext_1;
      entryValids_2 <= entryValidsNext_2;
      entryValids_3 <= entryValidsNext_3;
      if(logCondition) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // IssueQueueComponent.scala:L247
          `else
            if(!1'b0) begin
              $display("NOTE(IssueQueueComponent.scala:247):  [normal] LsuEU_IQ-3: STATUS - ValidCount=%x, allocateIn(valid=%x, ready=%x), issueOut(valid=%x, ready=%x)", currentValidCount, io_allocateIn_valid, io_allocateIn_ready, io_issueOut_valid, io_issueOut_ready); // IssueQueueComponent.scala:L247
            end
          `endif
        `endif
      end
      if(when_IssueQueueComponent_l256) begin
        if(entryValids_0) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] LsuEU_IQ-3: (LAST CYCLE) ENTRY[0] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_0_robPtr, entries_0_physDest_idx, entries_0_useSrc1, entries_0_src1Tag, entries_0_src1Ready, entries_0_useSrc2, entries_0_src2Tag, entries_0_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_1) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] LsuEU_IQ-3: (LAST CYCLE) ENTRY[1] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_1_robPtr, entries_1_physDest_idx, entries_1_useSrc1, entries_1_src1Tag, entries_1_src1Ready, entries_1_useSrc2, entries_1_src2Tag, entries_1_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_2) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] LsuEU_IQ-3: (LAST CYCLE) ENTRY[2] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_2_robPtr, entries_2_physDest_idx, entries_2_useSrc1, entries_2_src1Tag, entries_2_src1Ready, entries_2_useSrc2, entries_2_src2Tag, entries_2_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_3) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] LsuEU_IQ-3: (LAST CYCLE) ENTRY[3] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_3_robPtr, entries_3_physDest_idx, entries_3_useSrc1, entries_3_src1Tag, entries_3_src1Ready, entries_3_useSrc2, entries_3_src2Tag, entries_3_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
      end
    end
  end

  always @(posedge clk) begin
    entries_0_robPtr <= entriesNext_0_robPtr;
    entries_0_physDest_idx <= entriesNext_0_physDest_idx;
    entries_0_physDestIsFpr <= entriesNext_0_physDestIsFpr;
    entries_0_writesToPhysReg <= entriesNext_0_writesToPhysReg;
    entries_0_useSrc1 <= entriesNext_0_useSrc1;
    entries_0_src1Data <= entriesNext_0_src1Data;
    entries_0_src1Tag <= entriesNext_0_src1Tag;
    entries_0_src1Ready <= entriesNext_0_src1Ready;
    entries_0_src1IsFpr <= entriesNext_0_src1IsFpr;
    entries_0_useSrc2 <= entriesNext_0_useSrc2;
    entries_0_src2Data <= entriesNext_0_src2Data;
    entries_0_src2Tag <= entriesNext_0_src2Tag;
    entries_0_src2Ready <= entriesNext_0_src2Ready;
    entries_0_src2IsFpr <= entriesNext_0_src2IsFpr;
    entries_0_memCtrl_size <= entriesNext_0_memCtrl_size;
    entries_0_memCtrl_isSignedLoad <= entriesNext_0_memCtrl_isSignedLoad;
    entries_0_memCtrl_isStore <= entriesNext_0_memCtrl_isStore;
    entries_0_memCtrl_isLoadLinked <= entriesNext_0_memCtrl_isLoadLinked;
    entries_0_memCtrl_isStoreCond <= entriesNext_0_memCtrl_isStoreCond;
    entries_0_memCtrl_atomicOp <= entriesNext_0_memCtrl_atomicOp;
    entries_0_memCtrl_isFence <= entriesNext_0_memCtrl_isFence;
    entries_0_memCtrl_fenceMode <= entriesNext_0_memCtrl_fenceMode;
    entries_0_memCtrl_isCacheOp <= entriesNext_0_memCtrl_isCacheOp;
    entries_0_memCtrl_cacheOpType <= entriesNext_0_memCtrl_cacheOpType;
    entries_0_memCtrl_isPrefetch <= entriesNext_0_memCtrl_isPrefetch;
    entries_0_imm <= entriesNext_0_imm;
    entries_0_usePc <= entriesNext_0_usePc;
    entries_0_pcData <= entriesNext_0_pcData;
    entries_1_robPtr <= entriesNext_1_robPtr;
    entries_1_physDest_idx <= entriesNext_1_physDest_idx;
    entries_1_physDestIsFpr <= entriesNext_1_physDestIsFpr;
    entries_1_writesToPhysReg <= entriesNext_1_writesToPhysReg;
    entries_1_useSrc1 <= entriesNext_1_useSrc1;
    entries_1_src1Data <= entriesNext_1_src1Data;
    entries_1_src1Tag <= entriesNext_1_src1Tag;
    entries_1_src1Ready <= entriesNext_1_src1Ready;
    entries_1_src1IsFpr <= entriesNext_1_src1IsFpr;
    entries_1_useSrc2 <= entriesNext_1_useSrc2;
    entries_1_src2Data <= entriesNext_1_src2Data;
    entries_1_src2Tag <= entriesNext_1_src2Tag;
    entries_1_src2Ready <= entriesNext_1_src2Ready;
    entries_1_src2IsFpr <= entriesNext_1_src2IsFpr;
    entries_1_memCtrl_size <= entriesNext_1_memCtrl_size;
    entries_1_memCtrl_isSignedLoad <= entriesNext_1_memCtrl_isSignedLoad;
    entries_1_memCtrl_isStore <= entriesNext_1_memCtrl_isStore;
    entries_1_memCtrl_isLoadLinked <= entriesNext_1_memCtrl_isLoadLinked;
    entries_1_memCtrl_isStoreCond <= entriesNext_1_memCtrl_isStoreCond;
    entries_1_memCtrl_atomicOp <= entriesNext_1_memCtrl_atomicOp;
    entries_1_memCtrl_isFence <= entriesNext_1_memCtrl_isFence;
    entries_1_memCtrl_fenceMode <= entriesNext_1_memCtrl_fenceMode;
    entries_1_memCtrl_isCacheOp <= entriesNext_1_memCtrl_isCacheOp;
    entries_1_memCtrl_cacheOpType <= entriesNext_1_memCtrl_cacheOpType;
    entries_1_memCtrl_isPrefetch <= entriesNext_1_memCtrl_isPrefetch;
    entries_1_imm <= entriesNext_1_imm;
    entries_1_usePc <= entriesNext_1_usePc;
    entries_1_pcData <= entriesNext_1_pcData;
    entries_2_robPtr <= entriesNext_2_robPtr;
    entries_2_physDest_idx <= entriesNext_2_physDest_idx;
    entries_2_physDestIsFpr <= entriesNext_2_physDestIsFpr;
    entries_2_writesToPhysReg <= entriesNext_2_writesToPhysReg;
    entries_2_useSrc1 <= entriesNext_2_useSrc1;
    entries_2_src1Data <= entriesNext_2_src1Data;
    entries_2_src1Tag <= entriesNext_2_src1Tag;
    entries_2_src1Ready <= entriesNext_2_src1Ready;
    entries_2_src1IsFpr <= entriesNext_2_src1IsFpr;
    entries_2_useSrc2 <= entriesNext_2_useSrc2;
    entries_2_src2Data <= entriesNext_2_src2Data;
    entries_2_src2Tag <= entriesNext_2_src2Tag;
    entries_2_src2Ready <= entriesNext_2_src2Ready;
    entries_2_src2IsFpr <= entriesNext_2_src2IsFpr;
    entries_2_memCtrl_size <= entriesNext_2_memCtrl_size;
    entries_2_memCtrl_isSignedLoad <= entriesNext_2_memCtrl_isSignedLoad;
    entries_2_memCtrl_isStore <= entriesNext_2_memCtrl_isStore;
    entries_2_memCtrl_isLoadLinked <= entriesNext_2_memCtrl_isLoadLinked;
    entries_2_memCtrl_isStoreCond <= entriesNext_2_memCtrl_isStoreCond;
    entries_2_memCtrl_atomicOp <= entriesNext_2_memCtrl_atomicOp;
    entries_2_memCtrl_isFence <= entriesNext_2_memCtrl_isFence;
    entries_2_memCtrl_fenceMode <= entriesNext_2_memCtrl_fenceMode;
    entries_2_memCtrl_isCacheOp <= entriesNext_2_memCtrl_isCacheOp;
    entries_2_memCtrl_cacheOpType <= entriesNext_2_memCtrl_cacheOpType;
    entries_2_memCtrl_isPrefetch <= entriesNext_2_memCtrl_isPrefetch;
    entries_2_imm <= entriesNext_2_imm;
    entries_2_usePc <= entriesNext_2_usePc;
    entries_2_pcData <= entriesNext_2_pcData;
    entries_3_robPtr <= entriesNext_3_robPtr;
    entries_3_physDest_idx <= entriesNext_3_physDest_idx;
    entries_3_physDestIsFpr <= entriesNext_3_physDestIsFpr;
    entries_3_writesToPhysReg <= entriesNext_3_writesToPhysReg;
    entries_3_useSrc1 <= entriesNext_3_useSrc1;
    entries_3_src1Data <= entriesNext_3_src1Data;
    entries_3_src1Tag <= entriesNext_3_src1Tag;
    entries_3_src1Ready <= entriesNext_3_src1Ready;
    entries_3_src1IsFpr <= entriesNext_3_src1IsFpr;
    entries_3_useSrc2 <= entriesNext_3_useSrc2;
    entries_3_src2Data <= entriesNext_3_src2Data;
    entries_3_src2Tag <= entriesNext_3_src2Tag;
    entries_3_src2Ready <= entriesNext_3_src2Ready;
    entries_3_src2IsFpr <= entriesNext_3_src2IsFpr;
    entries_3_memCtrl_size <= entriesNext_3_memCtrl_size;
    entries_3_memCtrl_isSignedLoad <= entriesNext_3_memCtrl_isSignedLoad;
    entries_3_memCtrl_isStore <= entriesNext_3_memCtrl_isStore;
    entries_3_memCtrl_isLoadLinked <= entriesNext_3_memCtrl_isLoadLinked;
    entries_3_memCtrl_isStoreCond <= entriesNext_3_memCtrl_isStoreCond;
    entries_3_memCtrl_atomicOp <= entriesNext_3_memCtrl_atomicOp;
    entries_3_memCtrl_isFence <= entriesNext_3_memCtrl_isFence;
    entries_3_memCtrl_fenceMode <= entriesNext_3_memCtrl_fenceMode;
    entries_3_memCtrl_isCacheOp <= entriesNext_3_memCtrl_isCacheOp;
    entries_3_memCtrl_cacheOpType <= entriesNext_3_memCtrl_cacheOpType;
    entries_3_memCtrl_isPrefetch <= entriesNext_3_memCtrl_isPrefetch;
    entries_3_imm <= entriesNext_3_imm;
    entries_3_usePc <= entriesNext_3_usePc;
    entries_3_pcData <= entriesNext_3_pcData;
  end


endmodule

module IssueQueueComponent_2 (
  input  wire          io_allocateIn_valid,
  output wire          io_allocateIn_ready,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_pc,
  input  wire          io_allocateIn_payload_uop_decoded_isValid,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_uopCode,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_exeUnit,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_isa,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archDest_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archDest_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_writeArchDestEn,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archSrc1_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archSrc1_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_useArchSrc1,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archSrc2_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archSrc2_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_useArchSrc2,
  input  wire          io_allocateIn_payload_uop_decoded_usePcForAddr,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_imm,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_immUsage,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isSub,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isAdd,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isSigned,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_aluCtrl_logicOp,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isRight,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_memCtrl_size,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isStore,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_memCtrl_atomicOp,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isFence,
  input  wire [7:0]    io_allocateIn_payload_uop_decoded_memCtrl_fenceMode,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_branchCtrl_condition,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isJump,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isLink,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_opType,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond,
  input  wire [13:0]   io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isWrite,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isRead,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isExchange,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc,
  input  wire [19:0]   io_allocateIn_payload_uop_decoded_sysCtrl_sysCode,
  input  wire          io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn,
  input  wire          io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_decodeExceptionCode,
  input  wire          io_allocateIn_payload_uop_decoded_hasDecodeException,
  input  wire          io_allocateIn_payload_uop_decoded_isMicrocode,
  input  wire [7:0]    io_allocateIn_payload_uop_decoded_microcodeEntry,
  input  wire          io_allocateIn_payload_uop_decoded_isSerializing,
  input  wire          io_allocateIn_payload_uop_decoded_isBranchOrJump,
  input  wire          io_allocateIn_payload_uop_decoded_branchPrediction_isTaken,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_branchPrediction_target,
  input  wire          io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physSrc1_idx,
  input  wire          io_allocateIn_payload_uop_rename_physSrc1IsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physSrc2_idx,
  input  wire          io_allocateIn_payload_uop_rename_physSrc2IsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physDest_idx,
  input  wire          io_allocateIn_payload_uop_rename_physDestIsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_oldPhysDest_idx,
  input  wire          io_allocateIn_payload_uop_rename_oldPhysDestIsFpr,
  input  wire          io_allocateIn_payload_uop_rename_allocatesPhysDest,
  input  wire          io_allocateIn_payload_uop_rename_writesToPhysReg,
  input  wire [3:0]    io_allocateIn_payload_uop_robPtr,
  input  wire [15:0]   io_allocateIn_payload_uop_uniqueId,
  input  wire          io_allocateIn_payload_uop_dispatched,
  input  wire          io_allocateIn_payload_uop_executed,
  input  wire          io_allocateIn_payload_uop_hasException,
  input  wire [7:0]    io_allocateIn_payload_uop_exceptionCode,
  input  wire          io_allocateIn_payload_src1InitialReady,
  input  wire          io_allocateIn_payload_src2InitialReady,
  output wire          io_issueOut_valid,
  input  wire          io_issueOut_ready,
  output wire [3:0]    io_issueOut_payload_robPtr,
  output wire [5:0]    io_issueOut_payload_physDest_idx,
  output wire          io_issueOut_payload_physDestIsFpr,
  output wire          io_issueOut_payload_writesToPhysReg,
  output wire          io_issueOut_payload_useSrc1,
  output wire [31:0]   io_issueOut_payload_src1Data,
  output wire [5:0]    io_issueOut_payload_src1Tag,
  output wire          io_issueOut_payload_src1Ready,
  output wire          io_issueOut_payload_src1IsFpr,
  output wire          io_issueOut_payload_useSrc2,
  output wire [31:0]   io_issueOut_payload_src2Data,
  output wire [5:0]    io_issueOut_payload_src2Tag,
  output wire          io_issueOut_payload_src2Ready,
  output wire          io_issueOut_payload_src2IsFpr,
  output wire [4:0]    io_issueOut_payload_branchCtrl_condition,
  output wire          io_issueOut_payload_branchCtrl_isJump,
  output wire          io_issueOut_payload_branchCtrl_isLink,
  output wire [4:0]    io_issueOut_payload_branchCtrl_linkReg_idx,
  output wire [1:0]    io_issueOut_payload_branchCtrl_linkReg_rtype,
  output wire          io_issueOut_payload_branchCtrl_isIndirect,
  output wire [2:0]    io_issueOut_payload_branchCtrl_laCfIdx,
  output wire [31:0]   io_issueOut_payload_imm,
  output wire [31:0]   io_issueOut_payload_pc,
  output wire          io_issueOut_payload_branchPrediction_isTaken,
  output wire [31:0]   io_issueOut_payload_branchPrediction_target,
  output wire          io_issueOut_payload_branchPrediction_wasPredicted,
  input  wire          io_wakeupIn_0_valid,
  input  wire [5:0]    io_wakeupIn_0_payload_physRegIdx,
  input  wire          io_wakeupIn_1_valid,
  input  wire [5:0]    io_wakeupIn_1_payload_physRegIdx,
  input  wire          io_wakeupIn_2_valid,
  input  wire [5:0]    io_wakeupIn_2_payload_physRegIdx,
  input  wire          io_wakeupIn_3_valid,
  input  wire [5:0]    io_wakeupIn_3_payload_physRegIdx,
  input  wire          io_wakeupIn_4_valid,
  input  wire [5:0]    io_wakeupIn_4_payload_physRegIdx,
  input  wire          io_flush,
  input  wire          clk,
  input  wire          reset
);
  localparam BaseUopCode_NOP = 5'd0;
  localparam BaseUopCode_ILLEGAL = 5'd1;
  localparam BaseUopCode_ALU = 5'd2;
  localparam BaseUopCode_SHIFT = 5'd3;
  localparam BaseUopCode_MUL = 5'd4;
  localparam BaseUopCode_DIV = 5'd5;
  localparam BaseUopCode_LOAD = 5'd6;
  localparam BaseUopCode_STORE = 5'd7;
  localparam BaseUopCode_ATOMIC = 5'd8;
  localparam BaseUopCode_MEM_BARRIER = 5'd9;
  localparam BaseUopCode_PREFETCH = 5'd10;
  localparam BaseUopCode_BRANCH = 5'd11;
  localparam BaseUopCode_JUMP_REG = 5'd12;
  localparam BaseUopCode_JUMP_IMM = 5'd13;
  localparam BaseUopCode_SYSTEM_OP = 5'd14;
  localparam BaseUopCode_CSR_ACCESS = 5'd15;
  localparam BaseUopCode_FPU_ALU = 5'd16;
  localparam BaseUopCode_FPU_CVT = 5'd17;
  localparam BaseUopCode_FPU_CMP = 5'd18;
  localparam BaseUopCode_FPU_SEL = 5'd19;
  localparam BaseUopCode_LA_BITMANIP = 5'd20;
  localparam BaseUopCode_LA_CACOP = 5'd21;
  localparam BaseUopCode_LA_TLB = 5'd22;
  localparam BaseUopCode_IDLE = 5'd23;
  localparam ExeUnitType_NONE = 4'd0;
  localparam ExeUnitType_ALU_INT = 4'd1;
  localparam ExeUnitType_MUL_INT = 4'd2;
  localparam ExeUnitType_DIV_INT = 4'd3;
  localparam ExeUnitType_MEM = 4'd4;
  localparam ExeUnitType_BRU = 4'd5;
  localparam ExeUnitType_CSR = 4'd6;
  localparam ExeUnitType_FPU_ADD_MUL_CVT_CMP = 4'd7;
  localparam ExeUnitType_FPU_DIV_SQRT = 4'd8;
  localparam IsaType_UNKNOWN = 2'd0;
  localparam IsaType_DEMO = 2'd1;
  localparam IsaType_RISCV = 2'd2;
  localparam IsaType_LOONGARCH = 2'd3;
  localparam ArchRegType_GPR = 2'd0;
  localparam ArchRegType_FPR = 2'd1;
  localparam ArchRegType_CSR = 2'd2;
  localparam ArchRegType_LA_CF = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;
  localparam BranchCondition_NUL = 5'd0;
  localparam BranchCondition_EQ = 5'd1;
  localparam BranchCondition_NE = 5'd2;
  localparam BranchCondition_LT = 5'd3;
  localparam BranchCondition_GE = 5'd4;
  localparam BranchCondition_LTU = 5'd5;
  localparam BranchCondition_GEU = 5'd6;
  localparam BranchCondition_EQZ = 5'd7;
  localparam BranchCondition_NEZ = 5'd8;
  localparam BranchCondition_LTZ = 5'd9;
  localparam BranchCondition_GEZ = 5'd10;
  localparam BranchCondition_GTZ = 5'd11;
  localparam BranchCondition_LEZ = 5'd12;
  localparam BranchCondition_F_EQ = 5'd13;
  localparam BranchCondition_F_NE = 5'd14;
  localparam BranchCondition_F_LT = 5'd15;
  localparam BranchCondition_F_LE = 5'd16;
  localparam BranchCondition_F_UN = 5'd17;
  localparam BranchCondition_LA_CF_TRUE = 5'd18;
  localparam BranchCondition_LA_CF_FALSE = 5'd19;
  localparam DecodeExCode_INVALID = 2'd0;
  localparam DecodeExCode_FETCH_ERROR = 2'd1;
  localparam DecodeExCode_DECODE_ERROR = 2'd2;
  localparam DecodeExCode_OK = 2'd3;

  wire       [3:0]    _zz_issueRequestMask_ohFirst_masked;
  reg        [4:0]    _zz__zz_io_issueOut_payload_branchCtrl_condition;
  reg        [1:0]    _zz__zz_io_issueOut_payload_branchCtrl_linkReg_rtype;
  reg        [3:0]    _zz_io_issueOut_payload_robPtr;
  reg        [5:0]    _zz_io_issueOut_payload_physDest_idx;
  reg                 _zz_io_issueOut_payload_physDestIsFpr;
  reg                 _zz_io_issueOut_payload_writesToPhysReg;
  reg                 _zz_io_issueOut_payload_useSrc1;
  reg        [31:0]   _zz_io_issueOut_payload_src1Data;
  reg        [5:0]    _zz_io_issueOut_payload_src1Tag;
  reg                 _zz_io_issueOut_payload_src1Ready;
  reg                 _zz_io_issueOut_payload_src1IsFpr;
  reg                 _zz_io_issueOut_payload_useSrc2;
  reg        [31:0]   _zz_io_issueOut_payload_src2Data;
  reg        [5:0]    _zz_io_issueOut_payload_src2Tag;
  reg                 _zz_io_issueOut_payload_src2Ready;
  reg                 _zz_io_issueOut_payload_src2IsFpr;
  reg                 _zz_io_issueOut_payload_branchCtrl_isJump;
  reg                 _zz_io_issueOut_payload_branchCtrl_isLink;
  reg        [4:0]    _zz_io_issueOut_payload_branchCtrl_linkReg_idx;
  reg                 _zz_io_issueOut_payload_branchCtrl_isIndirect;
  reg        [2:0]    _zz_io_issueOut_payload_branchCtrl_laCfIdx;
  reg        [31:0]   _zz_io_issueOut_payload_imm;
  reg        [31:0]   _zz_io_issueOut_payload_pc;
  reg                 _zz_io_issueOut_payload_branchPrediction_isTaken;
  reg        [31:0]   _zz_io_issueOut_payload_branchPrediction_target;
  reg                 _zz_io_issueOut_payload_branchPrediction_wasPredicted;
  wire       [3:0]    _zz_allocationMask_1;
  reg        [2:0]    _zz_currentValidCount_8;
  wire       [2:0]    _zz_currentValidCount_9;
  reg        [2:0]    _zz_currentValidCount_10;
  wire       [2:0]    _zz_currentValidCount_11;
  wire       [0:0]    _zz_currentValidCount_12;
  reg        [3:0]    entries_0_robPtr;
  reg        [5:0]    entries_0_physDest_idx;
  reg                 entries_0_physDestIsFpr;
  reg                 entries_0_writesToPhysReg;
  reg                 entries_0_useSrc1;
  reg        [31:0]   entries_0_src1Data;
  reg        [5:0]    entries_0_src1Tag;
  reg                 entries_0_src1Ready;
  reg                 entries_0_src1IsFpr;
  reg                 entries_0_useSrc2;
  reg        [31:0]   entries_0_src2Data;
  reg        [5:0]    entries_0_src2Tag;
  reg                 entries_0_src2Ready;
  reg                 entries_0_src2IsFpr;
  reg        [4:0]    entries_0_branchCtrl_condition;
  reg                 entries_0_branchCtrl_isJump;
  reg                 entries_0_branchCtrl_isLink;
  reg        [4:0]    entries_0_branchCtrl_linkReg_idx;
  reg        [1:0]    entries_0_branchCtrl_linkReg_rtype;
  reg                 entries_0_branchCtrl_isIndirect;
  reg        [2:0]    entries_0_branchCtrl_laCfIdx;
  reg        [31:0]   entries_0_imm;
  reg        [31:0]   entries_0_pc;
  reg                 entries_0_branchPrediction_isTaken;
  reg        [31:0]   entries_0_branchPrediction_target;
  reg                 entries_0_branchPrediction_wasPredicted;
  reg        [3:0]    entries_1_robPtr;
  reg        [5:0]    entries_1_physDest_idx;
  reg                 entries_1_physDestIsFpr;
  reg                 entries_1_writesToPhysReg;
  reg                 entries_1_useSrc1;
  reg        [31:0]   entries_1_src1Data;
  reg        [5:0]    entries_1_src1Tag;
  reg                 entries_1_src1Ready;
  reg                 entries_1_src1IsFpr;
  reg                 entries_1_useSrc2;
  reg        [31:0]   entries_1_src2Data;
  reg        [5:0]    entries_1_src2Tag;
  reg                 entries_1_src2Ready;
  reg                 entries_1_src2IsFpr;
  reg        [4:0]    entries_1_branchCtrl_condition;
  reg                 entries_1_branchCtrl_isJump;
  reg                 entries_1_branchCtrl_isLink;
  reg        [4:0]    entries_1_branchCtrl_linkReg_idx;
  reg        [1:0]    entries_1_branchCtrl_linkReg_rtype;
  reg                 entries_1_branchCtrl_isIndirect;
  reg        [2:0]    entries_1_branchCtrl_laCfIdx;
  reg        [31:0]   entries_1_imm;
  reg        [31:0]   entries_1_pc;
  reg                 entries_1_branchPrediction_isTaken;
  reg        [31:0]   entries_1_branchPrediction_target;
  reg                 entries_1_branchPrediction_wasPredicted;
  reg        [3:0]    entries_2_robPtr;
  reg        [5:0]    entries_2_physDest_idx;
  reg                 entries_2_physDestIsFpr;
  reg                 entries_2_writesToPhysReg;
  reg                 entries_2_useSrc1;
  reg        [31:0]   entries_2_src1Data;
  reg        [5:0]    entries_2_src1Tag;
  reg                 entries_2_src1Ready;
  reg                 entries_2_src1IsFpr;
  reg                 entries_2_useSrc2;
  reg        [31:0]   entries_2_src2Data;
  reg        [5:0]    entries_2_src2Tag;
  reg                 entries_2_src2Ready;
  reg                 entries_2_src2IsFpr;
  reg        [4:0]    entries_2_branchCtrl_condition;
  reg                 entries_2_branchCtrl_isJump;
  reg                 entries_2_branchCtrl_isLink;
  reg        [4:0]    entries_2_branchCtrl_linkReg_idx;
  reg        [1:0]    entries_2_branchCtrl_linkReg_rtype;
  reg                 entries_2_branchCtrl_isIndirect;
  reg        [2:0]    entries_2_branchCtrl_laCfIdx;
  reg        [31:0]   entries_2_imm;
  reg        [31:0]   entries_2_pc;
  reg                 entries_2_branchPrediction_isTaken;
  reg        [31:0]   entries_2_branchPrediction_target;
  reg                 entries_2_branchPrediction_wasPredicted;
  reg        [3:0]    entries_3_robPtr;
  reg        [5:0]    entries_3_physDest_idx;
  reg                 entries_3_physDestIsFpr;
  reg                 entries_3_writesToPhysReg;
  reg                 entries_3_useSrc1;
  reg        [31:0]   entries_3_src1Data;
  reg        [5:0]    entries_3_src1Tag;
  reg                 entries_3_src1Ready;
  reg                 entries_3_src1IsFpr;
  reg                 entries_3_useSrc2;
  reg        [31:0]   entries_3_src2Data;
  reg        [5:0]    entries_3_src2Tag;
  reg                 entries_3_src2Ready;
  reg                 entries_3_src2IsFpr;
  reg        [4:0]    entries_3_branchCtrl_condition;
  reg                 entries_3_branchCtrl_isJump;
  reg                 entries_3_branchCtrl_isLink;
  reg        [4:0]    entries_3_branchCtrl_linkReg_idx;
  reg        [1:0]    entries_3_branchCtrl_linkReg_rtype;
  reg                 entries_3_branchCtrl_isIndirect;
  reg        [2:0]    entries_3_branchCtrl_laCfIdx;
  reg        [31:0]   entries_3_imm;
  reg        [31:0]   entries_3_pc;
  reg                 entries_3_branchPrediction_isTaken;
  reg        [31:0]   entries_3_branchPrediction_target;
  reg                 entries_3_branchPrediction_wasPredicted;
  reg                 entryValids_0;
  reg                 entryValids_1;
  reg                 entryValids_2;
  reg                 entryValids_3;
  wire                io_issueOut_fire;
  wire                localWakeupValid;
  reg        [3:0]    wokeUpSrc1Mask;
  reg        [3:0]    wokeUpSrc2Mask;
  wire                _zz_when_IssueQueueComponent_l103;
  wire                _zz_when_IssueQueueComponent_l106;
  wire                when_IssueQueueComponent_l103;
  wire                when_IssueQueueComponent_l106;
  wire                when_IssueQueueComponent_l113;
  wire                when_IssueQueueComponent_l116;
  wire                when_IssueQueueComponent_l113_1;
  wire                when_IssueQueueComponent_l116_1;
  wire                when_IssueQueueComponent_l113_2;
  wire                when_IssueQueueComponent_l116_2;
  wire                when_IssueQueueComponent_l113_3;
  wire                when_IssueQueueComponent_l116_3;
  wire                when_IssueQueueComponent_l113_4;
  wire                when_IssueQueueComponent_l116_4;
  wire                _zz_when_IssueQueueComponent_l103_1;
  wire                _zz_when_IssueQueueComponent_l106_1;
  wire                when_IssueQueueComponent_l103_1;
  wire                when_IssueQueueComponent_l106_1;
  wire                when_IssueQueueComponent_l113_5;
  wire                when_IssueQueueComponent_l116_5;
  wire                when_IssueQueueComponent_l113_6;
  wire                when_IssueQueueComponent_l116_6;
  wire                when_IssueQueueComponent_l113_7;
  wire                when_IssueQueueComponent_l116_7;
  wire                when_IssueQueueComponent_l113_8;
  wire                when_IssueQueueComponent_l116_8;
  wire                when_IssueQueueComponent_l113_9;
  wire                when_IssueQueueComponent_l116_9;
  wire                _zz_when_IssueQueueComponent_l103_2;
  wire                _zz_when_IssueQueueComponent_l106_2;
  wire                when_IssueQueueComponent_l103_2;
  wire                when_IssueQueueComponent_l106_2;
  wire                when_IssueQueueComponent_l113_10;
  wire                when_IssueQueueComponent_l116_10;
  wire                when_IssueQueueComponent_l113_11;
  wire                when_IssueQueueComponent_l116_11;
  wire                when_IssueQueueComponent_l113_12;
  wire                when_IssueQueueComponent_l116_12;
  wire                when_IssueQueueComponent_l113_13;
  wire                when_IssueQueueComponent_l116_13;
  wire                when_IssueQueueComponent_l113_14;
  wire                when_IssueQueueComponent_l116_14;
  wire                _zz_when_IssueQueueComponent_l103_3;
  wire                _zz_when_IssueQueueComponent_l106_3;
  wire                when_IssueQueueComponent_l103_3;
  wire                when_IssueQueueComponent_l106_3;
  wire                when_IssueQueueComponent_l113_15;
  wire                when_IssueQueueComponent_l116_15;
  wire                when_IssueQueueComponent_l113_16;
  wire                when_IssueQueueComponent_l116_16;
  wire                when_IssueQueueComponent_l113_17;
  wire                when_IssueQueueComponent_l116_17;
  wire                when_IssueQueueComponent_l113_18;
  wire                when_IssueQueueComponent_l116_18;
  wire                when_IssueQueueComponent_l113_19;
  wire                when_IssueQueueComponent_l116_19;
  wire                entriesReadyToIssue_0;
  wire                entriesReadyToIssue_1;
  wire                entriesReadyToIssue_2;
  wire                entriesReadyToIssue_3;
  wire       [3:0]    issueRequestMask;
  wire       [3:0]    issueRequestMask_ohFirst_input;
  wire       [3:0]    issueRequestMask_ohFirst_masked;
  wire       [3:0]    issueRequestOh;
  wire                _zz_issueIdx;
  wire                _zz_issueIdx_1;
  wire                _zz_issueIdx_2;
  wire       [1:0]    issueIdx;
  wire       [4:0]    _zz_io_issueOut_payload_branchCtrl_condition;
  wire       [1:0]    _zz_io_issueOut_payload_branchCtrl_linkReg_rtype;
  wire       [3:0]    freeSlotsMask;
  wire                hasSpaceForNewEntry;
  reg        [3:0]    firedSlotMask;
  wire       [3:0]    _zz_allocationMask;
  wire       [3:0]    allocationMask;
  wire                _zz_allocateIdx;
  wire                _zz_allocateIdx_1;
  wire                _zz_allocateIdx_2;
  wire       [1:0]    allocateIdx;
  reg        [3:0]    entriesNext_0_robPtr;
  reg        [5:0]    entriesNext_0_physDest_idx;
  reg                 entriesNext_0_physDestIsFpr;
  reg                 entriesNext_0_writesToPhysReg;
  reg                 entriesNext_0_useSrc1;
  reg        [31:0]   entriesNext_0_src1Data;
  reg        [5:0]    entriesNext_0_src1Tag;
  reg                 entriesNext_0_src1Ready;
  reg                 entriesNext_0_src1IsFpr;
  reg                 entriesNext_0_useSrc2;
  reg        [31:0]   entriesNext_0_src2Data;
  reg        [5:0]    entriesNext_0_src2Tag;
  reg                 entriesNext_0_src2Ready;
  reg                 entriesNext_0_src2IsFpr;
  reg        [4:0]    entriesNext_0_branchCtrl_condition;
  reg                 entriesNext_0_branchCtrl_isJump;
  reg                 entriesNext_0_branchCtrl_isLink;
  reg        [4:0]    entriesNext_0_branchCtrl_linkReg_idx;
  reg        [1:0]    entriesNext_0_branchCtrl_linkReg_rtype;
  reg                 entriesNext_0_branchCtrl_isIndirect;
  reg        [2:0]    entriesNext_0_branchCtrl_laCfIdx;
  reg        [31:0]   entriesNext_0_imm;
  reg        [31:0]   entriesNext_0_pc;
  reg                 entriesNext_0_branchPrediction_isTaken;
  reg        [31:0]   entriesNext_0_branchPrediction_target;
  reg                 entriesNext_0_branchPrediction_wasPredicted;
  reg        [3:0]    entriesNext_1_robPtr;
  reg        [5:0]    entriesNext_1_physDest_idx;
  reg                 entriesNext_1_physDestIsFpr;
  reg                 entriesNext_1_writesToPhysReg;
  reg                 entriesNext_1_useSrc1;
  reg        [31:0]   entriesNext_1_src1Data;
  reg        [5:0]    entriesNext_1_src1Tag;
  reg                 entriesNext_1_src1Ready;
  reg                 entriesNext_1_src1IsFpr;
  reg                 entriesNext_1_useSrc2;
  reg        [31:0]   entriesNext_1_src2Data;
  reg        [5:0]    entriesNext_1_src2Tag;
  reg                 entriesNext_1_src2Ready;
  reg                 entriesNext_1_src2IsFpr;
  reg        [4:0]    entriesNext_1_branchCtrl_condition;
  reg                 entriesNext_1_branchCtrl_isJump;
  reg                 entriesNext_1_branchCtrl_isLink;
  reg        [4:0]    entriesNext_1_branchCtrl_linkReg_idx;
  reg        [1:0]    entriesNext_1_branchCtrl_linkReg_rtype;
  reg                 entriesNext_1_branchCtrl_isIndirect;
  reg        [2:0]    entriesNext_1_branchCtrl_laCfIdx;
  reg        [31:0]   entriesNext_1_imm;
  reg        [31:0]   entriesNext_1_pc;
  reg                 entriesNext_1_branchPrediction_isTaken;
  reg        [31:0]   entriesNext_1_branchPrediction_target;
  reg                 entriesNext_1_branchPrediction_wasPredicted;
  reg        [3:0]    entriesNext_2_robPtr;
  reg        [5:0]    entriesNext_2_physDest_idx;
  reg                 entriesNext_2_physDestIsFpr;
  reg                 entriesNext_2_writesToPhysReg;
  reg                 entriesNext_2_useSrc1;
  reg        [31:0]   entriesNext_2_src1Data;
  reg        [5:0]    entriesNext_2_src1Tag;
  reg                 entriesNext_2_src1Ready;
  reg                 entriesNext_2_src1IsFpr;
  reg                 entriesNext_2_useSrc2;
  reg        [31:0]   entriesNext_2_src2Data;
  reg        [5:0]    entriesNext_2_src2Tag;
  reg                 entriesNext_2_src2Ready;
  reg                 entriesNext_2_src2IsFpr;
  reg        [4:0]    entriesNext_2_branchCtrl_condition;
  reg                 entriesNext_2_branchCtrl_isJump;
  reg                 entriesNext_2_branchCtrl_isLink;
  reg        [4:0]    entriesNext_2_branchCtrl_linkReg_idx;
  reg        [1:0]    entriesNext_2_branchCtrl_linkReg_rtype;
  reg                 entriesNext_2_branchCtrl_isIndirect;
  reg        [2:0]    entriesNext_2_branchCtrl_laCfIdx;
  reg        [31:0]   entriesNext_2_imm;
  reg        [31:0]   entriesNext_2_pc;
  reg                 entriesNext_2_branchPrediction_isTaken;
  reg        [31:0]   entriesNext_2_branchPrediction_target;
  reg                 entriesNext_2_branchPrediction_wasPredicted;
  reg        [3:0]    entriesNext_3_robPtr;
  reg        [5:0]    entriesNext_3_physDest_idx;
  reg                 entriesNext_3_physDestIsFpr;
  reg                 entriesNext_3_writesToPhysReg;
  reg                 entriesNext_3_useSrc1;
  reg        [31:0]   entriesNext_3_src1Data;
  reg        [5:0]    entriesNext_3_src1Tag;
  reg                 entriesNext_3_src1Ready;
  reg                 entriesNext_3_src1IsFpr;
  reg                 entriesNext_3_useSrc2;
  reg        [31:0]   entriesNext_3_src2Data;
  reg        [5:0]    entriesNext_3_src2Tag;
  reg                 entriesNext_3_src2Ready;
  reg                 entriesNext_3_src2IsFpr;
  reg        [4:0]    entriesNext_3_branchCtrl_condition;
  reg                 entriesNext_3_branchCtrl_isJump;
  reg                 entriesNext_3_branchCtrl_isLink;
  reg        [4:0]    entriesNext_3_branchCtrl_linkReg_idx;
  reg        [1:0]    entriesNext_3_branchCtrl_linkReg_rtype;
  reg                 entriesNext_3_branchCtrl_isIndirect;
  reg        [2:0]    entriesNext_3_branchCtrl_laCfIdx;
  reg        [31:0]   entriesNext_3_imm;
  reg        [31:0]   entriesNext_3_pc;
  reg                 entriesNext_3_branchPrediction_isTaken;
  reg        [31:0]   entriesNext_3_branchPrediction_target;
  reg                 entriesNext_3_branchPrediction_wasPredicted;
  reg                 entryValidsNext_0;
  reg                 entryValidsNext_1;
  reg                 entryValidsNext_2;
  reg                 entryValidsNext_3;
  wire                when_IssueQueueComponent_l186;
  wire                when_IssueQueueComponent_l187;
  wire                when_IssueQueueComponent_l186_1;
  wire                when_IssueQueueComponent_l187_1;
  wire                when_IssueQueueComponent_l186_2;
  wire                when_IssueQueueComponent_l187_2;
  wire                when_IssueQueueComponent_l186_3;
  wire                when_IssueQueueComponent_l187_3;
  wire       [3:0]    _zz_1;
  wire                io_allocateIn_fire;
  wire       [3:0]    _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_entriesNext_0_src1Ready;
  wire                _zz_entriesNext_0_src2Ready;
  wire       [3:0]    _zz_7;
  wire                when_IssueQueueComponent_l212;
  wire                when_IssueQueueComponent_l215;
  wire                when_IssueQueueComponent_l212_1;
  wire                when_IssueQueueComponent_l215_1;
  wire                when_IssueQueueComponent_l212_2;
  wire                when_IssueQueueComponent_l215_2;
  wire                when_IssueQueueComponent_l212_3;
  wire                when_IssueQueueComponent_l215_3;
  wire                when_IssueQueueComponent_l212_4;
  wire                when_IssueQueueComponent_l215_4;
  wire       [2:0]    _zz_currentValidCount;
  wire       [2:0]    _zz_currentValidCount_1;
  wire       [2:0]    _zz_currentValidCount_2;
  wire       [2:0]    _zz_currentValidCount_3;
  wire       [2:0]    _zz_currentValidCount_4;
  wire       [2:0]    _zz_currentValidCount_5;
  wire       [2:0]    _zz_currentValidCount_6;
  wire       [2:0]    _zz_currentValidCount_7;
  wire       [2:0]    currentValidCount;
  wire                logCondition;
  wire                when_IssueQueueComponent_l256;
  `ifndef SYNTHESIS
  reg [87:0] io_allocateIn_payload_uop_decoded_uopCode_string;
  reg [151:0] io_allocateIn_payload_uop_decoded_exeUnit_string;
  reg [71:0] io_allocateIn_payload_uop_decoded_isa_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] io_allocateIn_payload_uop_decoded_immUsage_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] io_allocateIn_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_allocateIn_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] io_issueOut_payload_branchCtrl_condition_string;
  reg [39:0] io_issueOut_payload_branchCtrl_linkReg_rtype_string;
  reg [87:0] entries_0_branchCtrl_condition_string;
  reg [39:0] entries_0_branchCtrl_linkReg_rtype_string;
  reg [87:0] entries_1_branchCtrl_condition_string;
  reg [39:0] entries_1_branchCtrl_linkReg_rtype_string;
  reg [87:0] entries_2_branchCtrl_condition_string;
  reg [39:0] entries_2_branchCtrl_linkReg_rtype_string;
  reg [87:0] entries_3_branchCtrl_condition_string;
  reg [39:0] entries_3_branchCtrl_linkReg_rtype_string;
  reg [87:0] _zz_io_issueOut_payload_branchCtrl_condition_string;
  reg [39:0] _zz_io_issueOut_payload_branchCtrl_linkReg_rtype_string;
  reg [87:0] entriesNext_0_branchCtrl_condition_string;
  reg [39:0] entriesNext_0_branchCtrl_linkReg_rtype_string;
  reg [87:0] entriesNext_1_branchCtrl_condition_string;
  reg [39:0] entriesNext_1_branchCtrl_linkReg_rtype_string;
  reg [87:0] entriesNext_2_branchCtrl_condition_string;
  reg [39:0] entriesNext_2_branchCtrl_linkReg_rtype_string;
  reg [87:0] entriesNext_3_branchCtrl_condition_string;
  reg [39:0] entriesNext_3_branchCtrl_linkReg_rtype_string;
  `endif


  assign _zz_issueRequestMask_ohFirst_masked = (issueRequestMask_ohFirst_input - 4'b0001);
  assign _zz_allocationMask_1 = (_zz_allocationMask - 4'b0001);
  assign _zz_currentValidCount_12 = entryValids_3;
  assign _zz_currentValidCount_11 = {2'd0, _zz_currentValidCount_12};
  assign _zz_currentValidCount_9 = {entryValids_2,{entryValids_1,entryValids_0}};
  always @(*) begin
    case(issueIdx)
      2'b00 : begin
        _zz__zz_io_issueOut_payload_branchCtrl_condition = entries_0_branchCtrl_condition;
        _zz__zz_io_issueOut_payload_branchCtrl_linkReg_rtype = entries_0_branchCtrl_linkReg_rtype;
        _zz_io_issueOut_payload_robPtr = entries_0_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_0_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_0_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_0_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_0_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_0_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_0_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_0_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_0_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_0_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_0_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_0_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_0_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_0_src2IsFpr;
        _zz_io_issueOut_payload_branchCtrl_isJump = entries_0_branchCtrl_isJump;
        _zz_io_issueOut_payload_branchCtrl_isLink = entries_0_branchCtrl_isLink;
        _zz_io_issueOut_payload_branchCtrl_linkReg_idx = entries_0_branchCtrl_linkReg_idx;
        _zz_io_issueOut_payload_branchCtrl_isIndirect = entries_0_branchCtrl_isIndirect;
        _zz_io_issueOut_payload_branchCtrl_laCfIdx = entries_0_branchCtrl_laCfIdx;
        _zz_io_issueOut_payload_imm = entries_0_imm;
        _zz_io_issueOut_payload_pc = entries_0_pc;
        _zz_io_issueOut_payload_branchPrediction_isTaken = entries_0_branchPrediction_isTaken;
        _zz_io_issueOut_payload_branchPrediction_target = entries_0_branchPrediction_target;
        _zz_io_issueOut_payload_branchPrediction_wasPredicted = entries_0_branchPrediction_wasPredicted;
      end
      2'b01 : begin
        _zz__zz_io_issueOut_payload_branchCtrl_condition = entries_1_branchCtrl_condition;
        _zz__zz_io_issueOut_payload_branchCtrl_linkReg_rtype = entries_1_branchCtrl_linkReg_rtype;
        _zz_io_issueOut_payload_robPtr = entries_1_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_1_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_1_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_1_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_1_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_1_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_1_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_1_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_1_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_1_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_1_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_1_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_1_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_1_src2IsFpr;
        _zz_io_issueOut_payload_branchCtrl_isJump = entries_1_branchCtrl_isJump;
        _zz_io_issueOut_payload_branchCtrl_isLink = entries_1_branchCtrl_isLink;
        _zz_io_issueOut_payload_branchCtrl_linkReg_idx = entries_1_branchCtrl_linkReg_idx;
        _zz_io_issueOut_payload_branchCtrl_isIndirect = entries_1_branchCtrl_isIndirect;
        _zz_io_issueOut_payload_branchCtrl_laCfIdx = entries_1_branchCtrl_laCfIdx;
        _zz_io_issueOut_payload_imm = entries_1_imm;
        _zz_io_issueOut_payload_pc = entries_1_pc;
        _zz_io_issueOut_payload_branchPrediction_isTaken = entries_1_branchPrediction_isTaken;
        _zz_io_issueOut_payload_branchPrediction_target = entries_1_branchPrediction_target;
        _zz_io_issueOut_payload_branchPrediction_wasPredicted = entries_1_branchPrediction_wasPredicted;
      end
      2'b10 : begin
        _zz__zz_io_issueOut_payload_branchCtrl_condition = entries_2_branchCtrl_condition;
        _zz__zz_io_issueOut_payload_branchCtrl_linkReg_rtype = entries_2_branchCtrl_linkReg_rtype;
        _zz_io_issueOut_payload_robPtr = entries_2_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_2_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_2_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_2_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_2_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_2_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_2_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_2_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_2_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_2_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_2_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_2_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_2_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_2_src2IsFpr;
        _zz_io_issueOut_payload_branchCtrl_isJump = entries_2_branchCtrl_isJump;
        _zz_io_issueOut_payload_branchCtrl_isLink = entries_2_branchCtrl_isLink;
        _zz_io_issueOut_payload_branchCtrl_linkReg_idx = entries_2_branchCtrl_linkReg_idx;
        _zz_io_issueOut_payload_branchCtrl_isIndirect = entries_2_branchCtrl_isIndirect;
        _zz_io_issueOut_payload_branchCtrl_laCfIdx = entries_2_branchCtrl_laCfIdx;
        _zz_io_issueOut_payload_imm = entries_2_imm;
        _zz_io_issueOut_payload_pc = entries_2_pc;
        _zz_io_issueOut_payload_branchPrediction_isTaken = entries_2_branchPrediction_isTaken;
        _zz_io_issueOut_payload_branchPrediction_target = entries_2_branchPrediction_target;
        _zz_io_issueOut_payload_branchPrediction_wasPredicted = entries_2_branchPrediction_wasPredicted;
      end
      default : begin
        _zz__zz_io_issueOut_payload_branchCtrl_condition = entries_3_branchCtrl_condition;
        _zz__zz_io_issueOut_payload_branchCtrl_linkReg_rtype = entries_3_branchCtrl_linkReg_rtype;
        _zz_io_issueOut_payload_robPtr = entries_3_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_3_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_3_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_3_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_3_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_3_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_3_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_3_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_3_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_3_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_3_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_3_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_3_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_3_src2IsFpr;
        _zz_io_issueOut_payload_branchCtrl_isJump = entries_3_branchCtrl_isJump;
        _zz_io_issueOut_payload_branchCtrl_isLink = entries_3_branchCtrl_isLink;
        _zz_io_issueOut_payload_branchCtrl_linkReg_idx = entries_3_branchCtrl_linkReg_idx;
        _zz_io_issueOut_payload_branchCtrl_isIndirect = entries_3_branchCtrl_isIndirect;
        _zz_io_issueOut_payload_branchCtrl_laCfIdx = entries_3_branchCtrl_laCfIdx;
        _zz_io_issueOut_payload_imm = entries_3_imm;
        _zz_io_issueOut_payload_pc = entries_3_pc;
        _zz_io_issueOut_payload_branchPrediction_isTaken = entries_3_branchPrediction_isTaken;
        _zz_io_issueOut_payload_branchPrediction_target = entries_3_branchPrediction_target;
        _zz_io_issueOut_payload_branchPrediction_wasPredicted = entries_3_branchPrediction_wasPredicted;
      end
    endcase
  end

  always @(*) begin
    case(_zz_currentValidCount_9)
      3'b000 : _zz_currentValidCount_8 = _zz_currentValidCount;
      3'b001 : _zz_currentValidCount_8 = _zz_currentValidCount_1;
      3'b010 : _zz_currentValidCount_8 = _zz_currentValidCount_2;
      3'b011 : _zz_currentValidCount_8 = _zz_currentValidCount_3;
      3'b100 : _zz_currentValidCount_8 = _zz_currentValidCount_4;
      3'b101 : _zz_currentValidCount_8 = _zz_currentValidCount_5;
      3'b110 : _zz_currentValidCount_8 = _zz_currentValidCount_6;
      default : _zz_currentValidCount_8 = _zz_currentValidCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_currentValidCount_11)
      3'b000 : _zz_currentValidCount_10 = _zz_currentValidCount;
      3'b001 : _zz_currentValidCount_10 = _zz_currentValidCount_1;
      3'b010 : _zz_currentValidCount_10 = _zz_currentValidCount_2;
      3'b011 : _zz_currentValidCount_10 = _zz_currentValidCount_3;
      3'b100 : _zz_currentValidCount_10 = _zz_currentValidCount_4;
      3'b101 : _zz_currentValidCount_10 = _zz_currentValidCount_5;
      3'b110 : _zz_currentValidCount_10 = _zz_currentValidCount_6;
      default : _zz_currentValidCount_10 = _zz_currentValidCount_7;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : io_allocateIn_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_allocateIn_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_allocateIn_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_allocateIn_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_allocateIn_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_allocateIn_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_allocateIn_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_allocateIn_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_allocateIn_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_allocateIn_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_allocateIn_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_allocateIn_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_allocateIn_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_allocateIn_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_allocateIn_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_allocateIn_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_allocateIn_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : io_allocateIn_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : io_allocateIn_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_allocateIn_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_allocateIn_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_allocateIn_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_allocateIn_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_allocateIn_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_allocateIn_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_isa)
      IsaType_UNKNOWN : io_allocateIn_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_allocateIn_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : io_allocateIn_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_allocateIn_payload_uop_decoded_isa_string = "LOONGARCH";
      default : io_allocateIn_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : io_allocateIn_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : io_allocateIn_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "D";
      default : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_branchCtrl_condition)
      BranchCondition_NUL : io_issueOut_payload_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_issueOut_payload_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_issueOut_payload_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_issueOut_payload_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_issueOut_payload_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_issueOut_payload_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_issueOut_payload_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_issueOut_payload_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_issueOut_payload_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_issueOut_payload_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_issueOut_payload_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_issueOut_payload_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_issueOut_payload_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_issueOut_payload_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_issueOut_payload_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_issueOut_payload_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_issueOut_payload_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_issueOut_payload_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_issueOut_payload_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_issueOut_payload_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_issueOut_payload_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_issueOut_payload_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_issueOut_payload_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_issueOut_payload_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_issueOut_payload_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_issueOut_payload_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_0_branchCtrl_condition)
      BranchCondition_NUL : entries_0_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entries_0_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entries_0_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entries_0_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entries_0_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entries_0_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entries_0_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entries_0_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entries_0_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entries_0_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entries_0_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entries_0_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entries_0_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entries_0_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entries_0_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entries_0_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entries_0_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entries_0_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entries_0_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entries_0_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entries_0_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_0_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entries_0_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_0_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_0_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_0_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entries_0_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_1_branchCtrl_condition)
      BranchCondition_NUL : entries_1_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entries_1_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entries_1_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entries_1_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entries_1_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entries_1_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entries_1_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entries_1_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entries_1_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entries_1_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entries_1_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entries_1_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entries_1_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entries_1_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entries_1_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entries_1_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entries_1_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entries_1_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entries_1_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entries_1_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entries_1_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_1_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entries_1_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_1_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_1_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_1_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entries_1_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_2_branchCtrl_condition)
      BranchCondition_NUL : entries_2_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entries_2_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entries_2_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entries_2_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entries_2_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entries_2_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entries_2_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entries_2_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entries_2_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entries_2_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entries_2_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entries_2_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entries_2_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entries_2_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entries_2_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entries_2_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entries_2_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entries_2_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entries_2_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entries_2_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entries_2_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_2_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entries_2_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_2_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_2_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_2_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entries_2_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_3_branchCtrl_condition)
      BranchCondition_NUL : entries_3_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entries_3_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entries_3_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entries_3_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entries_3_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entries_3_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entries_3_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entries_3_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entries_3_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entries_3_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entries_3_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entries_3_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entries_3_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entries_3_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entries_3_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entries_3_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entries_3_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entries_3_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entries_3_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entries_3_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entries_3_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_3_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entries_3_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_3_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_3_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_3_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entries_3_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_branchCtrl_condition)
      BranchCondition_NUL : _zz_io_issueOut_payload_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : _zz_io_issueOut_payload_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : _zz_io_issueOut_payload_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : _zz_io_issueOut_payload_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : _zz_io_issueOut_payload_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : _zz_io_issueOut_payload_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : _zz_io_issueOut_payload_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : _zz_io_issueOut_payload_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : _zz_io_issueOut_payload_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : _zz_io_issueOut_payload_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : _zz_io_issueOut_payload_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : _zz_io_issueOut_payload_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : _zz_io_issueOut_payload_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_io_issueOut_payload_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_io_issueOut_payload_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : _zz_io_issueOut_payload_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : _zz_io_issueOut_payload_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : _zz_io_issueOut_payload_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_io_issueOut_payload_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_io_issueOut_payload_branchCtrl_condition_string = "LA_CF_FALSE";
      default : _zz_io_issueOut_payload_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : _zz_io_issueOut_payload_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_issueOut_payload_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_issueOut_payload_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_issueOut_payload_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : _zz_io_issueOut_payload_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_branchCtrl_condition)
      BranchCondition_NUL : entriesNext_0_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entriesNext_0_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entriesNext_0_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entriesNext_0_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entriesNext_0_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entriesNext_0_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entriesNext_0_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entriesNext_0_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entriesNext_0_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entriesNext_0_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entriesNext_0_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entriesNext_0_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entriesNext_0_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entriesNext_0_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entriesNext_0_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entriesNext_0_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entriesNext_0_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entriesNext_0_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entriesNext_0_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entriesNext_0_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entriesNext_0_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entriesNext_0_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_0_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_0_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_0_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entriesNext_0_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_branchCtrl_condition)
      BranchCondition_NUL : entriesNext_1_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entriesNext_1_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entriesNext_1_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entriesNext_1_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entriesNext_1_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entriesNext_1_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entriesNext_1_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entriesNext_1_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entriesNext_1_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entriesNext_1_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entriesNext_1_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entriesNext_1_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entriesNext_1_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entriesNext_1_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entriesNext_1_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entriesNext_1_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entriesNext_1_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entriesNext_1_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entriesNext_1_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entriesNext_1_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entriesNext_1_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entriesNext_1_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_1_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_1_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_1_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entriesNext_1_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_branchCtrl_condition)
      BranchCondition_NUL : entriesNext_2_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entriesNext_2_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entriesNext_2_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entriesNext_2_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entriesNext_2_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entriesNext_2_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entriesNext_2_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entriesNext_2_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entriesNext_2_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entriesNext_2_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entriesNext_2_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entriesNext_2_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entriesNext_2_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entriesNext_2_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entriesNext_2_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entriesNext_2_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entriesNext_2_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entriesNext_2_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entriesNext_2_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entriesNext_2_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entriesNext_2_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entriesNext_2_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_2_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_2_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_2_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entriesNext_2_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_branchCtrl_condition)
      BranchCondition_NUL : entriesNext_3_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entriesNext_3_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entriesNext_3_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entriesNext_3_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entriesNext_3_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entriesNext_3_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entriesNext_3_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entriesNext_3_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entriesNext_3_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entriesNext_3_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entriesNext_3_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entriesNext_3_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entriesNext_3_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entriesNext_3_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entriesNext_3_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entriesNext_3_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entriesNext_3_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entriesNext_3_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entriesNext_3_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entriesNext_3_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entriesNext_3_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entriesNext_3_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_3_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_3_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_3_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entriesNext_3_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  `endif

  assign io_issueOut_fire = (io_issueOut_valid && io_issueOut_ready);
  assign localWakeupValid = (io_issueOut_fire && io_issueOut_payload_writesToPhysReg);
  always @(*) begin
    wokeUpSrc1Mask = 4'b0000;
    if(entryValids_0) begin
      if(when_IssueQueueComponent_l103) begin
        wokeUpSrc1Mask[0] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_1) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_2) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_3) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_4) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
    end
    if(entryValids_1) begin
      if(when_IssueQueueComponent_l103_1) begin
        wokeUpSrc1Mask[1] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_5) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_6) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_7) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_8) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_9) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
    end
    if(entryValids_2) begin
      if(when_IssueQueueComponent_l103_2) begin
        wokeUpSrc1Mask[2] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_10) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_11) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_12) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_13) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_14) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
    end
    if(entryValids_3) begin
      if(when_IssueQueueComponent_l103_3) begin
        wokeUpSrc1Mask[3] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_15) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_16) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_17) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_18) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_19) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    wokeUpSrc2Mask = 4'b0000;
    if(entryValids_0) begin
      if(when_IssueQueueComponent_l106) begin
        wokeUpSrc2Mask[0] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_1) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_2) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_3) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_4) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
    end
    if(entryValids_1) begin
      if(when_IssueQueueComponent_l106_1) begin
        wokeUpSrc2Mask[1] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_5) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_6) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_7) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_8) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_9) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
    end
    if(entryValids_2) begin
      if(when_IssueQueueComponent_l106_2) begin
        wokeUpSrc2Mask[2] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_10) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_11) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_12) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_13) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_14) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
    end
    if(entryValids_3) begin
      if(when_IssueQueueComponent_l106_3) begin
        wokeUpSrc2Mask[3] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_15) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_16) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_17) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_18) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_19) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
    end
  end

  assign _zz_when_IssueQueueComponent_l103 = ((! entries_0_src1Ready) && entries_0_useSrc1);
  assign _zz_when_IssueQueueComponent_l106 = ((! entries_0_src2Ready) && entries_0_useSrc2);
  assign when_IssueQueueComponent_l103 = ((_zz_when_IssueQueueComponent_l103 && localWakeupValid) && (entries_0_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106 = ((_zz_when_IssueQueueComponent_l106 && localWakeupValid) && (entries_0_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_1 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_1 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_2 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_2 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_3 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_3 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_4 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_4 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_1 = ((! entries_1_src1Ready) && entries_1_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_1 = ((! entries_1_src2Ready) && entries_1_useSrc2);
  assign when_IssueQueueComponent_l103_1 = ((_zz_when_IssueQueueComponent_l103_1 && localWakeupValid) && (entries_1_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_1 = ((_zz_when_IssueQueueComponent_l106_1 && localWakeupValid) && (entries_1_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_5 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_5 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_6 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_6 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_7 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_7 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_8 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_8 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_9 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_9 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_2 = ((! entries_2_src1Ready) && entries_2_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_2 = ((! entries_2_src2Ready) && entries_2_useSrc2);
  assign when_IssueQueueComponent_l103_2 = ((_zz_when_IssueQueueComponent_l103_2 && localWakeupValid) && (entries_2_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_2 = ((_zz_when_IssueQueueComponent_l106_2 && localWakeupValid) && (entries_2_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_10 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_10 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_11 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_11 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_12 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_12 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_13 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_13 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_14 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_14 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_3 = ((! entries_3_src1Ready) && entries_3_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_3 = ((! entries_3_src2Ready) && entries_3_useSrc2);
  assign when_IssueQueueComponent_l103_3 = ((_zz_when_IssueQueueComponent_l103_3 && localWakeupValid) && (entries_3_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_3 = ((_zz_when_IssueQueueComponent_l106_3 && localWakeupValid) && (entries_3_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_15 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_15 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_16 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_16 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_17 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_17 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_18 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_18 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_19 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_19 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign entriesReadyToIssue_0 = ((entryValids_0 && ((! entries_0_useSrc1) || entries_0_src1Ready)) && ((! entries_0_useSrc2) || entries_0_src2Ready));
  assign entriesReadyToIssue_1 = ((entryValids_1 && ((! entries_1_useSrc1) || entries_1_src1Ready)) && ((! entries_1_useSrc2) || entries_1_src2Ready));
  assign entriesReadyToIssue_2 = ((entryValids_2 && ((! entries_2_useSrc1) || entries_2_src1Ready)) && ((! entries_2_useSrc2) || entries_2_src2Ready));
  assign entriesReadyToIssue_3 = ((entryValids_3 && ((! entries_3_useSrc1) || entries_3_src1Ready)) && ((! entries_3_useSrc2) || entries_3_src2Ready));
  assign issueRequestMask = {entriesReadyToIssue_3,{entriesReadyToIssue_2,{entriesReadyToIssue_1,entriesReadyToIssue_0}}};
  assign issueRequestMask_ohFirst_input = issueRequestMask;
  assign issueRequestMask_ohFirst_masked = (issueRequestMask_ohFirst_input & (~ _zz_issueRequestMask_ohFirst_masked));
  assign issueRequestOh = issueRequestMask_ohFirst_masked;
  assign _zz_issueIdx = issueRequestOh[3];
  assign _zz_issueIdx_1 = (issueRequestOh[1] || _zz_issueIdx);
  assign _zz_issueIdx_2 = (issueRequestOh[2] || _zz_issueIdx);
  assign issueIdx = {_zz_issueIdx_2,_zz_issueIdx_1};
  assign io_issueOut_valid = ((|issueRequestOh) && (! io_flush));
  assign _zz_io_issueOut_payload_branchCtrl_condition = _zz__zz_io_issueOut_payload_branchCtrl_condition;
  assign _zz_io_issueOut_payload_branchCtrl_linkReg_rtype = _zz__zz_io_issueOut_payload_branchCtrl_linkReg_rtype;
  assign io_issueOut_payload_robPtr = _zz_io_issueOut_payload_robPtr;
  assign io_issueOut_payload_physDest_idx = _zz_io_issueOut_payload_physDest_idx;
  assign io_issueOut_payload_physDestIsFpr = _zz_io_issueOut_payload_physDestIsFpr;
  assign io_issueOut_payload_writesToPhysReg = _zz_io_issueOut_payload_writesToPhysReg;
  assign io_issueOut_payload_useSrc1 = _zz_io_issueOut_payload_useSrc1;
  assign io_issueOut_payload_src1Data = _zz_io_issueOut_payload_src1Data;
  assign io_issueOut_payload_src1Tag = _zz_io_issueOut_payload_src1Tag;
  assign io_issueOut_payload_src1Ready = _zz_io_issueOut_payload_src1Ready;
  assign io_issueOut_payload_src1IsFpr = _zz_io_issueOut_payload_src1IsFpr;
  assign io_issueOut_payload_useSrc2 = _zz_io_issueOut_payload_useSrc2;
  assign io_issueOut_payload_src2Data = _zz_io_issueOut_payload_src2Data;
  assign io_issueOut_payload_src2Tag = _zz_io_issueOut_payload_src2Tag;
  assign io_issueOut_payload_src2Ready = _zz_io_issueOut_payload_src2Ready;
  assign io_issueOut_payload_src2IsFpr = _zz_io_issueOut_payload_src2IsFpr;
  assign io_issueOut_payload_branchCtrl_condition = _zz_io_issueOut_payload_branchCtrl_condition;
  assign io_issueOut_payload_branchCtrl_isJump = _zz_io_issueOut_payload_branchCtrl_isJump;
  assign io_issueOut_payload_branchCtrl_isLink = _zz_io_issueOut_payload_branchCtrl_isLink;
  assign io_issueOut_payload_branchCtrl_linkReg_idx = _zz_io_issueOut_payload_branchCtrl_linkReg_idx;
  assign io_issueOut_payload_branchCtrl_linkReg_rtype = _zz_io_issueOut_payload_branchCtrl_linkReg_rtype;
  assign io_issueOut_payload_branchCtrl_isIndirect = _zz_io_issueOut_payload_branchCtrl_isIndirect;
  assign io_issueOut_payload_branchCtrl_laCfIdx = _zz_io_issueOut_payload_branchCtrl_laCfIdx;
  assign io_issueOut_payload_imm = _zz_io_issueOut_payload_imm;
  assign io_issueOut_payload_pc = _zz_io_issueOut_payload_pc;
  assign io_issueOut_payload_branchPrediction_isTaken = _zz_io_issueOut_payload_branchPrediction_isTaken;
  assign io_issueOut_payload_branchPrediction_target = _zz_io_issueOut_payload_branchPrediction_target;
  assign io_issueOut_payload_branchPrediction_wasPredicted = _zz_io_issueOut_payload_branchPrediction_wasPredicted;
  assign freeSlotsMask = {(! entryValids_3),{(! entryValids_2),{(! entryValids_1),(! entryValids_0)}}};
  assign hasSpaceForNewEntry = ((|freeSlotsMask) || io_issueOut_fire);
  assign io_allocateIn_ready = (hasSpaceForNewEntry && (! io_flush));
  always @(*) begin
    firedSlotMask = 4'b0000;
    if(io_issueOut_fire) begin
      firedSlotMask[issueIdx] = 1'b1;
    end
  end

  assign _zz_allocationMask = (freeSlotsMask | firedSlotMask);
  assign allocationMask = (_zz_allocationMask & (~ _zz_allocationMask_1));
  assign _zz_allocateIdx = allocationMask[3];
  assign _zz_allocateIdx_1 = (allocationMask[1] || _zz_allocateIdx);
  assign _zz_allocateIdx_2 = (allocationMask[2] || _zz_allocateIdx);
  assign allocateIdx = {_zz_allocateIdx_2,_zz_allocateIdx_1};
  always @(*) begin
    entriesNext_0_robPtr = entries_0_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_physDest_idx = entries_0_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_physDestIsFpr = entries_0_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_writesToPhysReg = entries_0_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_0_useSrc1 = entries_0_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Data = entries_0_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Tag = entries_0_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Ready = entries_0_src1Ready;
    if(when_IssueQueueComponent_l186) begin
      entriesNext_0_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_3) begin
        entriesNext_0_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1IsFpr = entries_0_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_useSrc2 = entries_0_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Data = entries_0_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Tag = entries_0_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Ready = entries_0_src2Ready;
    if(when_IssueQueueComponent_l187) begin
      entriesNext_0_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_3) begin
        entriesNext_0_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2IsFpr = entries_0_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchCtrl_condition = entries_0_branchCtrl_condition;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchCtrl_condition = io_allocateIn_payload_uop_decoded_branchCtrl_condition;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchCtrl_isJump = entries_0_branchCtrl_isJump;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchCtrl_isJump = io_allocateIn_payload_uop_decoded_branchCtrl_isJump;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchCtrl_isLink = entries_0_branchCtrl_isLink;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchCtrl_isLink = io_allocateIn_payload_uop_decoded_branchCtrl_isLink;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchCtrl_linkReg_idx = entries_0_branchCtrl_linkReg_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchCtrl_linkReg_idx = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchCtrl_linkReg_rtype = entries_0_branchCtrl_linkReg_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchCtrl_linkReg_rtype = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchCtrl_isIndirect = entries_0_branchCtrl_isIndirect;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchCtrl_isIndirect = io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchCtrl_laCfIdx = entries_0_branchCtrl_laCfIdx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchCtrl_laCfIdx = io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_imm = entries_0_imm;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_0_pc = entries_0_pc;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_pc = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchPrediction_isTaken = entries_0_branchPrediction_isTaken;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchPrediction_isTaken = io_allocateIn_payload_uop_decoded_branchPrediction_isTaken;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchPrediction_target = entries_0_branchPrediction_target;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchPrediction_target = io_allocateIn_payload_uop_decoded_branchPrediction_target;
      end
    end
  end

  always @(*) begin
    entriesNext_0_branchPrediction_wasPredicted = entries_0_branchPrediction_wasPredicted;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_branchPrediction_wasPredicted = io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted;
      end
    end
  end

  always @(*) begin
    entriesNext_1_robPtr = entries_1_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_physDest_idx = entries_1_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_physDestIsFpr = entries_1_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_writesToPhysReg = entries_1_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_1_useSrc1 = entries_1_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Data = entries_1_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Tag = entries_1_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Ready = entries_1_src1Ready;
    if(when_IssueQueueComponent_l186_1) begin
      entriesNext_1_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_4) begin
        entriesNext_1_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1IsFpr = entries_1_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_useSrc2 = entries_1_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Data = entries_1_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Tag = entries_1_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Ready = entries_1_src2Ready;
    if(when_IssueQueueComponent_l187_1) begin
      entriesNext_1_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_4) begin
        entriesNext_1_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2IsFpr = entries_1_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchCtrl_condition = entries_1_branchCtrl_condition;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchCtrl_condition = io_allocateIn_payload_uop_decoded_branchCtrl_condition;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchCtrl_isJump = entries_1_branchCtrl_isJump;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchCtrl_isJump = io_allocateIn_payload_uop_decoded_branchCtrl_isJump;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchCtrl_isLink = entries_1_branchCtrl_isLink;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchCtrl_isLink = io_allocateIn_payload_uop_decoded_branchCtrl_isLink;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchCtrl_linkReg_idx = entries_1_branchCtrl_linkReg_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchCtrl_linkReg_idx = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchCtrl_linkReg_rtype = entries_1_branchCtrl_linkReg_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchCtrl_linkReg_rtype = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchCtrl_isIndirect = entries_1_branchCtrl_isIndirect;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchCtrl_isIndirect = io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchCtrl_laCfIdx = entries_1_branchCtrl_laCfIdx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchCtrl_laCfIdx = io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_imm = entries_1_imm;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_1_pc = entries_1_pc;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_pc = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchPrediction_isTaken = entries_1_branchPrediction_isTaken;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchPrediction_isTaken = io_allocateIn_payload_uop_decoded_branchPrediction_isTaken;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchPrediction_target = entries_1_branchPrediction_target;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchPrediction_target = io_allocateIn_payload_uop_decoded_branchPrediction_target;
      end
    end
  end

  always @(*) begin
    entriesNext_1_branchPrediction_wasPredicted = entries_1_branchPrediction_wasPredicted;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_branchPrediction_wasPredicted = io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted;
      end
    end
  end

  always @(*) begin
    entriesNext_2_robPtr = entries_2_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_physDest_idx = entries_2_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_physDestIsFpr = entries_2_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_writesToPhysReg = entries_2_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_2_useSrc1 = entries_2_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Data = entries_2_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Tag = entries_2_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Ready = entries_2_src1Ready;
    if(when_IssueQueueComponent_l186_2) begin
      entriesNext_2_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_5) begin
        entriesNext_2_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1IsFpr = entries_2_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_useSrc2 = entries_2_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Data = entries_2_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Tag = entries_2_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Ready = entries_2_src2Ready;
    if(when_IssueQueueComponent_l187_2) begin
      entriesNext_2_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_5) begin
        entriesNext_2_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2IsFpr = entries_2_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchCtrl_condition = entries_2_branchCtrl_condition;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchCtrl_condition = io_allocateIn_payload_uop_decoded_branchCtrl_condition;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchCtrl_isJump = entries_2_branchCtrl_isJump;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchCtrl_isJump = io_allocateIn_payload_uop_decoded_branchCtrl_isJump;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchCtrl_isLink = entries_2_branchCtrl_isLink;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchCtrl_isLink = io_allocateIn_payload_uop_decoded_branchCtrl_isLink;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchCtrl_linkReg_idx = entries_2_branchCtrl_linkReg_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchCtrl_linkReg_idx = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchCtrl_linkReg_rtype = entries_2_branchCtrl_linkReg_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchCtrl_linkReg_rtype = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchCtrl_isIndirect = entries_2_branchCtrl_isIndirect;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchCtrl_isIndirect = io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchCtrl_laCfIdx = entries_2_branchCtrl_laCfIdx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchCtrl_laCfIdx = io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_imm = entries_2_imm;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_2_pc = entries_2_pc;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_pc = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchPrediction_isTaken = entries_2_branchPrediction_isTaken;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchPrediction_isTaken = io_allocateIn_payload_uop_decoded_branchPrediction_isTaken;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchPrediction_target = entries_2_branchPrediction_target;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchPrediction_target = io_allocateIn_payload_uop_decoded_branchPrediction_target;
      end
    end
  end

  always @(*) begin
    entriesNext_2_branchPrediction_wasPredicted = entries_2_branchPrediction_wasPredicted;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_branchPrediction_wasPredicted = io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted;
      end
    end
  end

  always @(*) begin
    entriesNext_3_robPtr = entries_3_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_physDest_idx = entries_3_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_physDestIsFpr = entries_3_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_writesToPhysReg = entries_3_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_3_useSrc1 = entries_3_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Data = entries_3_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Tag = entries_3_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Ready = entries_3_src1Ready;
    if(when_IssueQueueComponent_l186_3) begin
      entriesNext_3_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_6) begin
        entriesNext_3_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1IsFpr = entries_3_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_useSrc2 = entries_3_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Data = entries_3_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Tag = entries_3_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Ready = entries_3_src2Ready;
    if(when_IssueQueueComponent_l187_3) begin
      entriesNext_3_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_6) begin
        entriesNext_3_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2IsFpr = entries_3_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchCtrl_condition = entries_3_branchCtrl_condition;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchCtrl_condition = io_allocateIn_payload_uop_decoded_branchCtrl_condition;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchCtrl_isJump = entries_3_branchCtrl_isJump;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchCtrl_isJump = io_allocateIn_payload_uop_decoded_branchCtrl_isJump;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchCtrl_isLink = entries_3_branchCtrl_isLink;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchCtrl_isLink = io_allocateIn_payload_uop_decoded_branchCtrl_isLink;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchCtrl_linkReg_idx = entries_3_branchCtrl_linkReg_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchCtrl_linkReg_idx = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchCtrl_linkReg_rtype = entries_3_branchCtrl_linkReg_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchCtrl_linkReg_rtype = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchCtrl_isIndirect = entries_3_branchCtrl_isIndirect;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchCtrl_isIndirect = io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchCtrl_laCfIdx = entries_3_branchCtrl_laCfIdx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchCtrl_laCfIdx = io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_imm = entries_3_imm;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_3_pc = entries_3_pc;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_pc = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchPrediction_isTaken = entries_3_branchPrediction_isTaken;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchPrediction_isTaken = io_allocateIn_payload_uop_decoded_branchPrediction_isTaken;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchPrediction_target = entries_3_branchPrediction_target;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchPrediction_target = io_allocateIn_payload_uop_decoded_branchPrediction_target;
      end
    end
  end

  always @(*) begin
    entriesNext_3_branchPrediction_wasPredicted = entries_3_branchPrediction_wasPredicted;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_branchPrediction_wasPredicted = io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted;
      end
    end
  end

  always @(*) begin
    entryValidsNext_0 = entryValids_0;
    if(io_issueOut_fire) begin
      if(_zz_1[0]) begin
        entryValidsNext_0 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[0]) begin
        entryValidsNext_0 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_0 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_1 = entryValids_1;
    if(io_issueOut_fire) begin
      if(_zz_1[1]) begin
        entryValidsNext_1 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[1]) begin
        entryValidsNext_1 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_1 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_2 = entryValids_2;
    if(io_issueOut_fire) begin
      if(_zz_1[2]) begin
        entryValidsNext_2 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[2]) begin
        entryValidsNext_2 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_2 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_3 = entryValids_3;
    if(io_issueOut_fire) begin
      if(_zz_1[3]) begin
        entryValidsNext_3 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[3]) begin
        entryValidsNext_3 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_3 = 1'b0;
    end
  end

  assign when_IssueQueueComponent_l186 = wokeUpSrc1Mask[0];
  assign when_IssueQueueComponent_l187 = wokeUpSrc2Mask[0];
  assign when_IssueQueueComponent_l186_1 = wokeUpSrc1Mask[1];
  assign when_IssueQueueComponent_l187_1 = wokeUpSrc2Mask[1];
  assign when_IssueQueueComponent_l186_2 = wokeUpSrc1Mask[2];
  assign when_IssueQueueComponent_l187_2 = wokeUpSrc2Mask[2];
  assign when_IssueQueueComponent_l186_3 = wokeUpSrc1Mask[3];
  assign when_IssueQueueComponent_l187_3 = wokeUpSrc2Mask[3];
  assign _zz_1 = ({3'd0,1'b1} <<< issueIdx);
  assign io_allocateIn_fire = (io_allocateIn_valid && io_allocateIn_ready);
  assign _zz_2 = ({3'd0,1'b1} <<< allocateIdx);
  assign _zz_3 = _zz_2[0];
  assign _zz_4 = _zz_2[1];
  assign _zz_5 = _zz_2[2];
  assign _zz_6 = _zz_2[3];
  assign _zz_entriesNext_0_src1Ready = (! io_allocateIn_payload_uop_decoded_useArchSrc1);
  assign _zz_entriesNext_0_src2Ready = (! io_allocateIn_payload_uop_decoded_useArchSrc2);
  assign _zz_7 = ({3'd0,1'b1} <<< allocateIdx);
  assign when_IssueQueueComponent_l212 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l215 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_1 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_1 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_2 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_2 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_3 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_3 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_4 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_4 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_currentValidCount = 3'b000;
  assign _zz_currentValidCount_1 = 3'b001;
  assign _zz_currentValidCount_2 = 3'b001;
  assign _zz_currentValidCount_3 = 3'b010;
  assign _zz_currentValidCount_4 = 3'b001;
  assign _zz_currentValidCount_5 = 3'b010;
  assign _zz_currentValidCount_6 = 3'b010;
  assign _zz_currentValidCount_7 = 3'b011;
  assign currentValidCount = (_zz_currentValidCount_8 + _zz_currentValidCount_10);
  assign logCondition = (io_allocateIn_fire || io_issueOut_fire);
  assign when_IssueQueueComponent_l256 = (logCondition && (3'b000 < currentValidCount));
  always @(posedge clk) begin
    if(reset) begin
      entryValids_0 <= 1'b0;
      entryValids_1 <= 1'b0;
      entryValids_2 <= 1'b0;
      entryValids_3 <= 1'b0;
    end else begin
      entryValids_0 <= entryValidsNext_0;
      entryValids_1 <= entryValidsNext_1;
      entryValids_2 <= entryValidsNext_2;
      entryValids_3 <= entryValidsNext_3;
      if(logCondition) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // IssueQueueComponent.scala:L247
          `else
            if(!1'b0) begin
              $display("NOTE(IssueQueueComponent.scala:247):  [normal] BranchEU_IQ-2: STATUS - ValidCount=%x, allocateIn(valid=%x, ready=%x), issueOut(valid=%x, ready=%x)", currentValidCount, io_allocateIn_valid, io_allocateIn_ready, io_issueOut_valid, io_issueOut_ready); // IssueQueueComponent.scala:L247
            end
          `endif
        `endif
      end
      if(when_IssueQueueComponent_l256) begin
        if(entryValids_0) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] BranchEU_IQ-2: (LAST CYCLE) ENTRY[0] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_0_robPtr, entries_0_physDest_idx, entries_0_useSrc1, entries_0_src1Tag, entries_0_src1Ready, entries_0_useSrc2, entries_0_src2Tag, entries_0_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_1) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] BranchEU_IQ-2: (LAST CYCLE) ENTRY[1] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_1_robPtr, entries_1_physDest_idx, entries_1_useSrc1, entries_1_src1Tag, entries_1_src1Ready, entries_1_useSrc2, entries_1_src2Tag, entries_1_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_2) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] BranchEU_IQ-2: (LAST CYCLE) ENTRY[2] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_2_robPtr, entries_2_physDest_idx, entries_2_useSrc1, entries_2_src1Tag, entries_2_src1Ready, entries_2_useSrc2, entries_2_src2Tag, entries_2_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_3) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] BranchEU_IQ-2: (LAST CYCLE) ENTRY[3] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_3_robPtr, entries_3_physDest_idx, entries_3_useSrc1, entries_3_src1Tag, entries_3_src1Ready, entries_3_useSrc2, entries_3_src2Tag, entries_3_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
      end
    end
  end

  always @(posedge clk) begin
    entries_0_robPtr <= entriesNext_0_robPtr;
    entries_0_physDest_idx <= entriesNext_0_physDest_idx;
    entries_0_physDestIsFpr <= entriesNext_0_physDestIsFpr;
    entries_0_writesToPhysReg <= entriesNext_0_writesToPhysReg;
    entries_0_useSrc1 <= entriesNext_0_useSrc1;
    entries_0_src1Data <= entriesNext_0_src1Data;
    entries_0_src1Tag <= entriesNext_0_src1Tag;
    entries_0_src1Ready <= entriesNext_0_src1Ready;
    entries_0_src1IsFpr <= entriesNext_0_src1IsFpr;
    entries_0_useSrc2 <= entriesNext_0_useSrc2;
    entries_0_src2Data <= entriesNext_0_src2Data;
    entries_0_src2Tag <= entriesNext_0_src2Tag;
    entries_0_src2Ready <= entriesNext_0_src2Ready;
    entries_0_src2IsFpr <= entriesNext_0_src2IsFpr;
    entries_0_branchCtrl_condition <= entriesNext_0_branchCtrl_condition;
    entries_0_branchCtrl_isJump <= entriesNext_0_branchCtrl_isJump;
    entries_0_branchCtrl_isLink <= entriesNext_0_branchCtrl_isLink;
    entries_0_branchCtrl_linkReg_idx <= entriesNext_0_branchCtrl_linkReg_idx;
    entries_0_branchCtrl_linkReg_rtype <= entriesNext_0_branchCtrl_linkReg_rtype;
    entries_0_branchCtrl_isIndirect <= entriesNext_0_branchCtrl_isIndirect;
    entries_0_branchCtrl_laCfIdx <= entriesNext_0_branchCtrl_laCfIdx;
    entries_0_imm <= entriesNext_0_imm;
    entries_0_pc <= entriesNext_0_pc;
    entries_0_branchPrediction_isTaken <= entriesNext_0_branchPrediction_isTaken;
    entries_0_branchPrediction_target <= entriesNext_0_branchPrediction_target;
    entries_0_branchPrediction_wasPredicted <= entriesNext_0_branchPrediction_wasPredicted;
    entries_1_robPtr <= entriesNext_1_robPtr;
    entries_1_physDest_idx <= entriesNext_1_physDest_idx;
    entries_1_physDestIsFpr <= entriesNext_1_physDestIsFpr;
    entries_1_writesToPhysReg <= entriesNext_1_writesToPhysReg;
    entries_1_useSrc1 <= entriesNext_1_useSrc1;
    entries_1_src1Data <= entriesNext_1_src1Data;
    entries_1_src1Tag <= entriesNext_1_src1Tag;
    entries_1_src1Ready <= entriesNext_1_src1Ready;
    entries_1_src1IsFpr <= entriesNext_1_src1IsFpr;
    entries_1_useSrc2 <= entriesNext_1_useSrc2;
    entries_1_src2Data <= entriesNext_1_src2Data;
    entries_1_src2Tag <= entriesNext_1_src2Tag;
    entries_1_src2Ready <= entriesNext_1_src2Ready;
    entries_1_src2IsFpr <= entriesNext_1_src2IsFpr;
    entries_1_branchCtrl_condition <= entriesNext_1_branchCtrl_condition;
    entries_1_branchCtrl_isJump <= entriesNext_1_branchCtrl_isJump;
    entries_1_branchCtrl_isLink <= entriesNext_1_branchCtrl_isLink;
    entries_1_branchCtrl_linkReg_idx <= entriesNext_1_branchCtrl_linkReg_idx;
    entries_1_branchCtrl_linkReg_rtype <= entriesNext_1_branchCtrl_linkReg_rtype;
    entries_1_branchCtrl_isIndirect <= entriesNext_1_branchCtrl_isIndirect;
    entries_1_branchCtrl_laCfIdx <= entriesNext_1_branchCtrl_laCfIdx;
    entries_1_imm <= entriesNext_1_imm;
    entries_1_pc <= entriesNext_1_pc;
    entries_1_branchPrediction_isTaken <= entriesNext_1_branchPrediction_isTaken;
    entries_1_branchPrediction_target <= entriesNext_1_branchPrediction_target;
    entries_1_branchPrediction_wasPredicted <= entriesNext_1_branchPrediction_wasPredicted;
    entries_2_robPtr <= entriesNext_2_robPtr;
    entries_2_physDest_idx <= entriesNext_2_physDest_idx;
    entries_2_physDestIsFpr <= entriesNext_2_physDestIsFpr;
    entries_2_writesToPhysReg <= entriesNext_2_writesToPhysReg;
    entries_2_useSrc1 <= entriesNext_2_useSrc1;
    entries_2_src1Data <= entriesNext_2_src1Data;
    entries_2_src1Tag <= entriesNext_2_src1Tag;
    entries_2_src1Ready <= entriesNext_2_src1Ready;
    entries_2_src1IsFpr <= entriesNext_2_src1IsFpr;
    entries_2_useSrc2 <= entriesNext_2_useSrc2;
    entries_2_src2Data <= entriesNext_2_src2Data;
    entries_2_src2Tag <= entriesNext_2_src2Tag;
    entries_2_src2Ready <= entriesNext_2_src2Ready;
    entries_2_src2IsFpr <= entriesNext_2_src2IsFpr;
    entries_2_branchCtrl_condition <= entriesNext_2_branchCtrl_condition;
    entries_2_branchCtrl_isJump <= entriesNext_2_branchCtrl_isJump;
    entries_2_branchCtrl_isLink <= entriesNext_2_branchCtrl_isLink;
    entries_2_branchCtrl_linkReg_idx <= entriesNext_2_branchCtrl_linkReg_idx;
    entries_2_branchCtrl_linkReg_rtype <= entriesNext_2_branchCtrl_linkReg_rtype;
    entries_2_branchCtrl_isIndirect <= entriesNext_2_branchCtrl_isIndirect;
    entries_2_branchCtrl_laCfIdx <= entriesNext_2_branchCtrl_laCfIdx;
    entries_2_imm <= entriesNext_2_imm;
    entries_2_pc <= entriesNext_2_pc;
    entries_2_branchPrediction_isTaken <= entriesNext_2_branchPrediction_isTaken;
    entries_2_branchPrediction_target <= entriesNext_2_branchPrediction_target;
    entries_2_branchPrediction_wasPredicted <= entriesNext_2_branchPrediction_wasPredicted;
    entries_3_robPtr <= entriesNext_3_robPtr;
    entries_3_physDest_idx <= entriesNext_3_physDest_idx;
    entries_3_physDestIsFpr <= entriesNext_3_physDestIsFpr;
    entries_3_writesToPhysReg <= entriesNext_3_writesToPhysReg;
    entries_3_useSrc1 <= entriesNext_3_useSrc1;
    entries_3_src1Data <= entriesNext_3_src1Data;
    entries_3_src1Tag <= entriesNext_3_src1Tag;
    entries_3_src1Ready <= entriesNext_3_src1Ready;
    entries_3_src1IsFpr <= entriesNext_3_src1IsFpr;
    entries_3_useSrc2 <= entriesNext_3_useSrc2;
    entries_3_src2Data <= entriesNext_3_src2Data;
    entries_3_src2Tag <= entriesNext_3_src2Tag;
    entries_3_src2Ready <= entriesNext_3_src2Ready;
    entries_3_src2IsFpr <= entriesNext_3_src2IsFpr;
    entries_3_branchCtrl_condition <= entriesNext_3_branchCtrl_condition;
    entries_3_branchCtrl_isJump <= entriesNext_3_branchCtrl_isJump;
    entries_3_branchCtrl_isLink <= entriesNext_3_branchCtrl_isLink;
    entries_3_branchCtrl_linkReg_idx <= entriesNext_3_branchCtrl_linkReg_idx;
    entries_3_branchCtrl_linkReg_rtype <= entriesNext_3_branchCtrl_linkReg_rtype;
    entries_3_branchCtrl_isIndirect <= entriesNext_3_branchCtrl_isIndirect;
    entries_3_branchCtrl_laCfIdx <= entriesNext_3_branchCtrl_laCfIdx;
    entries_3_imm <= entriesNext_3_imm;
    entries_3_pc <= entriesNext_3_pc;
    entries_3_branchPrediction_isTaken <= entriesNext_3_branchPrediction_isTaken;
    entries_3_branchPrediction_target <= entriesNext_3_branchPrediction_target;
    entries_3_branchPrediction_wasPredicted <= entriesNext_3_branchPrediction_wasPredicted;
  end


endmodule

module IssueQueueComponent_1 (
  input  wire          io_allocateIn_valid,
  output wire          io_allocateIn_ready,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_pc,
  input  wire          io_allocateIn_payload_uop_decoded_isValid,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_uopCode,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_exeUnit,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_isa,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archDest_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archDest_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_writeArchDestEn,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archSrc1_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archSrc1_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_useArchSrc1,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archSrc2_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archSrc2_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_useArchSrc2,
  input  wire          io_allocateIn_payload_uop_decoded_usePcForAddr,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_imm,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_immUsage,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isSub,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isAdd,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isSigned,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_aluCtrl_logicOp,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isRight,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_memCtrl_size,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isStore,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_memCtrl_atomicOp,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isFence,
  input  wire [7:0]    io_allocateIn_payload_uop_decoded_memCtrl_fenceMode,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_branchCtrl_condition,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isJump,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isLink,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_opType,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond,
  input  wire [13:0]   io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isWrite,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isRead,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isExchange,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc,
  input  wire [19:0]   io_allocateIn_payload_uop_decoded_sysCtrl_sysCode,
  input  wire          io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn,
  input  wire          io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_decodeExceptionCode,
  input  wire          io_allocateIn_payload_uop_decoded_hasDecodeException,
  input  wire          io_allocateIn_payload_uop_decoded_isMicrocode,
  input  wire [7:0]    io_allocateIn_payload_uop_decoded_microcodeEntry,
  input  wire          io_allocateIn_payload_uop_decoded_isSerializing,
  input  wire          io_allocateIn_payload_uop_decoded_isBranchOrJump,
  input  wire          io_allocateIn_payload_uop_decoded_branchPrediction_isTaken,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_branchPrediction_target,
  input  wire          io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physSrc1_idx,
  input  wire          io_allocateIn_payload_uop_rename_physSrc1IsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physSrc2_idx,
  input  wire          io_allocateIn_payload_uop_rename_physSrc2IsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physDest_idx,
  input  wire          io_allocateIn_payload_uop_rename_physDestIsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_oldPhysDest_idx,
  input  wire          io_allocateIn_payload_uop_rename_oldPhysDestIsFpr,
  input  wire          io_allocateIn_payload_uop_rename_allocatesPhysDest,
  input  wire          io_allocateIn_payload_uop_rename_writesToPhysReg,
  input  wire [3:0]    io_allocateIn_payload_uop_robPtr,
  input  wire [15:0]   io_allocateIn_payload_uop_uniqueId,
  input  wire          io_allocateIn_payload_uop_dispatched,
  input  wire          io_allocateIn_payload_uop_executed,
  input  wire          io_allocateIn_payload_uop_hasException,
  input  wire [7:0]    io_allocateIn_payload_uop_exceptionCode,
  input  wire          io_allocateIn_payload_src1InitialReady,
  input  wire          io_allocateIn_payload_src2InitialReady,
  output wire          io_issueOut_valid,
  input  wire          io_issueOut_ready,
  output wire [31:0]   io_issueOut_payload_uop_decoded_pc,
  output wire          io_issueOut_payload_uop_decoded_isValid,
  output wire [4:0]    io_issueOut_payload_uop_decoded_uopCode,
  output wire [3:0]    io_issueOut_payload_uop_decoded_exeUnit,
  output wire [1:0]    io_issueOut_payload_uop_decoded_isa,
  output wire [4:0]    io_issueOut_payload_uop_decoded_archDest_idx,
  output wire [1:0]    io_issueOut_payload_uop_decoded_archDest_rtype,
  output wire          io_issueOut_payload_uop_decoded_writeArchDestEn,
  output wire [4:0]    io_issueOut_payload_uop_decoded_archSrc1_idx,
  output wire [1:0]    io_issueOut_payload_uop_decoded_archSrc1_rtype,
  output wire          io_issueOut_payload_uop_decoded_useArchSrc1,
  output wire [4:0]    io_issueOut_payload_uop_decoded_archSrc2_idx,
  output wire [1:0]    io_issueOut_payload_uop_decoded_archSrc2_rtype,
  output wire          io_issueOut_payload_uop_decoded_useArchSrc2,
  output wire          io_issueOut_payload_uop_decoded_usePcForAddr,
  output wire [31:0]   io_issueOut_payload_uop_decoded_imm,
  output wire [2:0]    io_issueOut_payload_uop_decoded_immUsage,
  output wire          io_issueOut_payload_uop_decoded_aluCtrl_valid,
  output wire          io_issueOut_payload_uop_decoded_aluCtrl_isSub,
  output wire          io_issueOut_payload_uop_decoded_aluCtrl_isAdd,
  output wire          io_issueOut_payload_uop_decoded_aluCtrl_isSigned,
  output wire [1:0]    io_issueOut_payload_uop_decoded_aluCtrl_logicOp,
  output wire          io_issueOut_payload_uop_decoded_shiftCtrl_valid,
  output wire          io_issueOut_payload_uop_decoded_shiftCtrl_isRight,
  output wire          io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic,
  output wire          io_issueOut_payload_uop_decoded_shiftCtrl_isRotate,
  output wire          io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord,
  output wire          io_issueOut_payload_uop_decoded_mulDivCtrl_valid,
  output wire          io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv,
  output wire          io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned,
  output wire          io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp,
  output wire [1:0]    io_issueOut_payload_uop_decoded_memCtrl_size,
  output wire          io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad,
  output wire          io_issueOut_payload_uop_decoded_memCtrl_isStore,
  output wire          io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked,
  output wire          io_issueOut_payload_uop_decoded_memCtrl_isStoreCond,
  output wire [4:0]    io_issueOut_payload_uop_decoded_memCtrl_atomicOp,
  output wire          io_issueOut_payload_uop_decoded_memCtrl_isFence,
  output wire [7:0]    io_issueOut_payload_uop_decoded_memCtrl_fenceMode,
  output wire          io_issueOut_payload_uop_decoded_memCtrl_isCacheOp,
  output wire [4:0]    io_issueOut_payload_uop_decoded_memCtrl_cacheOpType,
  output wire          io_issueOut_payload_uop_decoded_memCtrl_isPrefetch,
  output wire [4:0]    io_issueOut_payload_uop_decoded_branchCtrl_condition,
  output wire          io_issueOut_payload_uop_decoded_branchCtrl_isJump,
  output wire          io_issueOut_payload_uop_decoded_branchCtrl_isLink,
  output wire [4:0]    io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx,
  output wire [1:0]    io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype,
  output wire          io_issueOut_payload_uop_decoded_branchCtrl_isIndirect,
  output wire [2:0]    io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx,
  output wire [3:0]    io_issueOut_payload_uop_decoded_fpuCtrl_opType,
  output wire [1:0]    io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1,
  output wire [1:0]    io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2,
  output wire [1:0]    io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest,
  output wire [2:0]    io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode,
  output wire          io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest,
  output wire          io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt,
  output wire          io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1,
  output wire [4:0]    io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond,
  output wire [13:0]   io_issueOut_payload_uop_decoded_csrCtrl_csrAddr,
  output wire          io_issueOut_payload_uop_decoded_csrCtrl_isWrite,
  output wire          io_issueOut_payload_uop_decoded_csrCtrl_isRead,
  output wire          io_issueOut_payload_uop_decoded_csrCtrl_isExchange,
  output wire          io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc,
  output wire [19:0]   io_issueOut_payload_uop_decoded_sysCtrl_sysCode,
  output wire          io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn,
  output wire          io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp,
  output wire [3:0]    io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType,
  output wire [1:0]    io_issueOut_payload_uop_decoded_decodeExceptionCode,
  output wire          io_issueOut_payload_uop_decoded_hasDecodeException,
  output wire          io_issueOut_payload_uop_decoded_isMicrocode,
  output wire [7:0]    io_issueOut_payload_uop_decoded_microcodeEntry,
  output wire          io_issueOut_payload_uop_decoded_isSerializing,
  output wire          io_issueOut_payload_uop_decoded_isBranchOrJump,
  output wire          io_issueOut_payload_uop_decoded_branchPrediction_isTaken,
  output wire [31:0]   io_issueOut_payload_uop_decoded_branchPrediction_target,
  output wire          io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted,
  output wire [5:0]    io_issueOut_payload_uop_rename_physSrc1_idx,
  output wire          io_issueOut_payload_uop_rename_physSrc1IsFpr,
  output wire [5:0]    io_issueOut_payload_uop_rename_physSrc2_idx,
  output wire          io_issueOut_payload_uop_rename_physSrc2IsFpr,
  output wire [5:0]    io_issueOut_payload_uop_rename_physDest_idx,
  output wire          io_issueOut_payload_uop_rename_physDestIsFpr,
  output wire [5:0]    io_issueOut_payload_uop_rename_oldPhysDest_idx,
  output wire          io_issueOut_payload_uop_rename_oldPhysDestIsFpr,
  output wire          io_issueOut_payload_uop_rename_allocatesPhysDest,
  output wire          io_issueOut_payload_uop_rename_writesToPhysReg,
  output wire [3:0]    io_issueOut_payload_uop_robPtr,
  output wire [15:0]   io_issueOut_payload_uop_uniqueId,
  output wire          io_issueOut_payload_uop_dispatched,
  output wire          io_issueOut_payload_uop_executed,
  output wire          io_issueOut_payload_uop_hasException,
  output wire [7:0]    io_issueOut_payload_uop_exceptionCode,
  output wire [3:0]    io_issueOut_payload_robPtr,
  output wire [5:0]    io_issueOut_payload_physDest_idx,
  output wire          io_issueOut_payload_physDestIsFpr,
  output wire          io_issueOut_payload_writesToPhysReg,
  output wire          io_issueOut_payload_useSrc1,
  output wire [31:0]   io_issueOut_payload_src1Data,
  output wire [5:0]    io_issueOut_payload_src1Tag,
  output wire          io_issueOut_payload_src1Ready,
  output wire          io_issueOut_payload_src1IsFpr,
  output wire          io_issueOut_payload_useSrc2,
  output wire [31:0]   io_issueOut_payload_src2Data,
  output wire [5:0]    io_issueOut_payload_src2Tag,
  output wire          io_issueOut_payload_src2Ready,
  output wire          io_issueOut_payload_src2IsFpr,
  output wire          io_issueOut_payload_mulDivCtrl_valid,
  output wire          io_issueOut_payload_mulDivCtrl_isDiv,
  output wire          io_issueOut_payload_mulDivCtrl_isSigned,
  output wire          io_issueOut_payload_mulDivCtrl_isWordOp,
  input  wire          io_wakeupIn_0_valid,
  input  wire [5:0]    io_wakeupIn_0_payload_physRegIdx,
  input  wire          io_wakeupIn_1_valid,
  input  wire [5:0]    io_wakeupIn_1_payload_physRegIdx,
  input  wire          io_wakeupIn_2_valid,
  input  wire [5:0]    io_wakeupIn_2_payload_physRegIdx,
  input  wire          io_wakeupIn_3_valid,
  input  wire [5:0]    io_wakeupIn_3_payload_physRegIdx,
  input  wire          io_wakeupIn_4_valid,
  input  wire [5:0]    io_wakeupIn_4_payload_physRegIdx,
  input  wire          io_flush,
  input  wire          clk,
  input  wire          reset
);
  localparam BaseUopCode_NOP = 5'd0;
  localparam BaseUopCode_ILLEGAL = 5'd1;
  localparam BaseUopCode_ALU = 5'd2;
  localparam BaseUopCode_SHIFT = 5'd3;
  localparam BaseUopCode_MUL = 5'd4;
  localparam BaseUopCode_DIV = 5'd5;
  localparam BaseUopCode_LOAD = 5'd6;
  localparam BaseUopCode_STORE = 5'd7;
  localparam BaseUopCode_ATOMIC = 5'd8;
  localparam BaseUopCode_MEM_BARRIER = 5'd9;
  localparam BaseUopCode_PREFETCH = 5'd10;
  localparam BaseUopCode_BRANCH = 5'd11;
  localparam BaseUopCode_JUMP_REG = 5'd12;
  localparam BaseUopCode_JUMP_IMM = 5'd13;
  localparam BaseUopCode_SYSTEM_OP = 5'd14;
  localparam BaseUopCode_CSR_ACCESS = 5'd15;
  localparam BaseUopCode_FPU_ALU = 5'd16;
  localparam BaseUopCode_FPU_CVT = 5'd17;
  localparam BaseUopCode_FPU_CMP = 5'd18;
  localparam BaseUopCode_FPU_SEL = 5'd19;
  localparam BaseUopCode_LA_BITMANIP = 5'd20;
  localparam BaseUopCode_LA_CACOP = 5'd21;
  localparam BaseUopCode_LA_TLB = 5'd22;
  localparam BaseUopCode_IDLE = 5'd23;
  localparam ExeUnitType_NONE = 4'd0;
  localparam ExeUnitType_ALU_INT = 4'd1;
  localparam ExeUnitType_MUL_INT = 4'd2;
  localparam ExeUnitType_DIV_INT = 4'd3;
  localparam ExeUnitType_MEM = 4'd4;
  localparam ExeUnitType_BRU = 4'd5;
  localparam ExeUnitType_CSR = 4'd6;
  localparam ExeUnitType_FPU_ADD_MUL_CVT_CMP = 4'd7;
  localparam ExeUnitType_FPU_DIV_SQRT = 4'd8;
  localparam IsaType_UNKNOWN = 2'd0;
  localparam IsaType_DEMO = 2'd1;
  localparam IsaType_RISCV = 2'd2;
  localparam IsaType_LOONGARCH = 2'd3;
  localparam ArchRegType_GPR = 2'd0;
  localparam ArchRegType_FPR = 2'd1;
  localparam ArchRegType_CSR = 2'd2;
  localparam ArchRegType_LA_CF = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;
  localparam BranchCondition_NUL = 5'd0;
  localparam BranchCondition_EQ = 5'd1;
  localparam BranchCondition_NE = 5'd2;
  localparam BranchCondition_LT = 5'd3;
  localparam BranchCondition_GE = 5'd4;
  localparam BranchCondition_LTU = 5'd5;
  localparam BranchCondition_GEU = 5'd6;
  localparam BranchCondition_EQZ = 5'd7;
  localparam BranchCondition_NEZ = 5'd8;
  localparam BranchCondition_LTZ = 5'd9;
  localparam BranchCondition_GEZ = 5'd10;
  localparam BranchCondition_GTZ = 5'd11;
  localparam BranchCondition_LEZ = 5'd12;
  localparam BranchCondition_F_EQ = 5'd13;
  localparam BranchCondition_F_NE = 5'd14;
  localparam BranchCondition_F_LT = 5'd15;
  localparam BranchCondition_F_LE = 5'd16;
  localparam BranchCondition_F_UN = 5'd17;
  localparam BranchCondition_LA_CF_TRUE = 5'd18;
  localparam BranchCondition_LA_CF_FALSE = 5'd19;
  localparam DecodeExCode_INVALID = 2'd0;
  localparam DecodeExCode_FETCH_ERROR = 2'd1;
  localparam DecodeExCode_DECODE_ERROR = 2'd2;
  localparam DecodeExCode_OK = 2'd3;

  wire       [3:0]    _zz_issueRequestMask_ohFirst_masked;
  reg        [4:0]    _zz__zz_io_issueOut_payload_uop_decoded_uopCode;
  reg        [3:0]    _zz__zz_io_issueOut_payload_uop_decoded_exeUnit;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_isa;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_archDest_rtype;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_archSrc1_rtype;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_archSrc2_rtype;
  reg        [2:0]    _zz__zz_io_issueOut_payload_uop_decoded_immUsage;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_memCtrl_size;
  reg        [4:0]    _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_condition;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [1:0]    _zz__zz_io_issueOut_payload_uop_decoded_decodeExceptionCode;
  reg        [31:0]   _zz_io_issueOut_payload_uop_decoded_pc;
  reg                 _zz_io_issueOut_payload_uop_decoded_isValid;
  reg        [4:0]    _zz_io_issueOut_payload_uop_decoded_archDest_idx;
  reg                 _zz_io_issueOut_payload_uop_decoded_writeArchDestEn;
  reg        [4:0]    _zz_io_issueOut_payload_uop_decoded_archSrc1_idx;
  reg                 _zz_io_issueOut_payload_uop_decoded_useArchSrc1;
  reg        [4:0]    _zz_io_issueOut_payload_uop_decoded_archSrc2_idx;
  reg                 _zz_io_issueOut_payload_uop_decoded_useArchSrc2;
  reg                 _zz_io_issueOut_payload_uop_decoded_usePcForAddr;
  reg        [31:0]   _zz_io_issueOut_payload_uop_decoded_imm;
  reg                 _zz_io_issueOut_payload_uop_decoded_aluCtrl_valid;
  reg                 _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSub;
  reg                 _zz_io_issueOut_payload_uop_decoded_aluCtrl_isAdd;
  reg                 _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSigned;
  reg                 _zz_io_issueOut_payload_uop_decoded_shiftCtrl_valid;
  reg                 _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRight;
  reg                 _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic;
  reg                 _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate;
  reg                 _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_valid;
  reg                 _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv;
  reg                 _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned;
  reg                 _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp;
  reg                 _zz_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad;
  reg                 _zz_io_issueOut_payload_uop_decoded_memCtrl_isStore;
  reg                 _zz_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked;
  reg                 _zz_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    _zz_io_issueOut_payload_uop_decoded_memCtrl_atomicOp;
  reg                 _zz_io_issueOut_payload_uop_decoded_memCtrl_isFence;
  reg        [7:0]    _zz_io_issueOut_payload_uop_decoded_memCtrl_fenceMode;
  reg                 _zz_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    _zz_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType;
  reg                 _zz_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch;
  reg                 _zz_io_issueOut_payload_uop_decoded_branchCtrl_isJump;
  reg                 _zz_io_issueOut_payload_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx;
  reg                 _zz_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    _zz_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    _zz_io_issueOut_payload_uop_decoded_fpuCtrl_opType;
  reg        [2:0]    _zz_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode;
  reg                 _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   _zz_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr;
  reg                 _zz_io_issueOut_payload_uop_decoded_csrCtrl_isWrite;
  reg                 _zz_io_issueOut_payload_uop_decoded_csrCtrl_isRead;
  reg                 _zz_io_issueOut_payload_uop_decoded_csrCtrl_isExchange;
  reg                 _zz_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   _zz_io_issueOut_payload_uop_decoded_sysCtrl_sysCode;
  reg                 _zz_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 _zz_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    _zz_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType;
  reg                 _zz_io_issueOut_payload_uop_decoded_hasDecodeException;
  reg                 _zz_io_issueOut_payload_uop_decoded_isMicrocode;
  reg        [7:0]    _zz_io_issueOut_payload_uop_decoded_microcodeEntry;
  reg                 _zz_io_issueOut_payload_uop_decoded_isSerializing;
  reg                 _zz_io_issueOut_payload_uop_decoded_isBranchOrJump;
  reg                 _zz_io_issueOut_payload_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   _zz_io_issueOut_payload_uop_decoded_branchPrediction_target;
  reg                 _zz_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    _zz_io_issueOut_payload_uop_rename_physSrc1_idx;
  reg                 _zz_io_issueOut_payload_uop_rename_physSrc1IsFpr;
  reg        [5:0]    _zz_io_issueOut_payload_uop_rename_physSrc2_idx;
  reg                 _zz_io_issueOut_payload_uop_rename_physSrc2IsFpr;
  reg        [5:0]    _zz_io_issueOut_payload_uop_rename_physDest_idx;
  reg                 _zz_io_issueOut_payload_uop_rename_physDestIsFpr;
  reg        [5:0]    _zz_io_issueOut_payload_uop_rename_oldPhysDest_idx;
  reg                 _zz_io_issueOut_payload_uop_rename_oldPhysDestIsFpr;
  reg                 _zz_io_issueOut_payload_uop_rename_allocatesPhysDest;
  reg                 _zz_io_issueOut_payload_uop_rename_writesToPhysReg;
  reg        [3:0]    _zz_io_issueOut_payload_uop_robPtr;
  reg        [15:0]   _zz_io_issueOut_payload_uop_uniqueId;
  reg                 _zz_io_issueOut_payload_uop_dispatched;
  reg                 _zz_io_issueOut_payload_uop_executed;
  reg                 _zz_io_issueOut_payload_uop_hasException;
  reg        [7:0]    _zz_io_issueOut_payload_uop_exceptionCode;
  reg        [3:0]    _zz_io_issueOut_payload_robPtr;
  reg        [5:0]    _zz_io_issueOut_payload_physDest_idx;
  reg                 _zz_io_issueOut_payload_physDestIsFpr;
  reg                 _zz_io_issueOut_payload_writesToPhysReg;
  reg                 _zz_io_issueOut_payload_useSrc1;
  reg        [31:0]   _zz_io_issueOut_payload_src1Data;
  reg        [5:0]    _zz_io_issueOut_payload_src1Tag;
  reg                 _zz_io_issueOut_payload_src1Ready;
  reg                 _zz_io_issueOut_payload_src1IsFpr;
  reg                 _zz_io_issueOut_payload_useSrc2;
  reg        [31:0]   _zz_io_issueOut_payload_src2Data;
  reg        [5:0]    _zz_io_issueOut_payload_src2Tag;
  reg                 _zz_io_issueOut_payload_src2Ready;
  reg                 _zz_io_issueOut_payload_src2IsFpr;
  reg                 _zz_io_issueOut_payload_mulDivCtrl_valid;
  reg                 _zz_io_issueOut_payload_mulDivCtrl_isDiv;
  reg                 _zz_io_issueOut_payload_mulDivCtrl_isSigned;
  reg                 _zz_io_issueOut_payload_mulDivCtrl_isWordOp;
  wire       [3:0]    _zz_allocationMask_1;
  reg        [2:0]    _zz_currentValidCount_8;
  wire       [2:0]    _zz_currentValidCount_9;
  reg        [2:0]    _zz_currentValidCount_10;
  wire       [2:0]    _zz_currentValidCount_11;
  wire       [0:0]    _zz_currentValidCount_12;
  reg        [31:0]   entries_0_uop_decoded_pc;
  reg                 entries_0_uop_decoded_isValid;
  reg        [4:0]    entries_0_uop_decoded_uopCode;
  reg        [3:0]    entries_0_uop_decoded_exeUnit;
  reg        [1:0]    entries_0_uop_decoded_isa;
  reg        [4:0]    entries_0_uop_decoded_archDest_idx;
  reg        [1:0]    entries_0_uop_decoded_archDest_rtype;
  reg                 entries_0_uop_decoded_writeArchDestEn;
  reg        [4:0]    entries_0_uop_decoded_archSrc1_idx;
  reg        [1:0]    entries_0_uop_decoded_archSrc1_rtype;
  reg                 entries_0_uop_decoded_useArchSrc1;
  reg        [4:0]    entries_0_uop_decoded_archSrc2_idx;
  reg        [1:0]    entries_0_uop_decoded_archSrc2_rtype;
  reg                 entries_0_uop_decoded_useArchSrc2;
  reg                 entries_0_uop_decoded_usePcForAddr;
  reg        [31:0]   entries_0_uop_decoded_imm;
  reg        [2:0]    entries_0_uop_decoded_immUsage;
  reg                 entries_0_uop_decoded_aluCtrl_valid;
  reg                 entries_0_uop_decoded_aluCtrl_isSub;
  reg                 entries_0_uop_decoded_aluCtrl_isAdd;
  reg                 entries_0_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    entries_0_uop_decoded_aluCtrl_logicOp;
  reg                 entries_0_uop_decoded_shiftCtrl_valid;
  reg                 entries_0_uop_decoded_shiftCtrl_isRight;
  reg                 entries_0_uop_decoded_shiftCtrl_isArithmetic;
  reg                 entries_0_uop_decoded_shiftCtrl_isRotate;
  reg                 entries_0_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 entries_0_uop_decoded_mulDivCtrl_valid;
  reg                 entries_0_uop_decoded_mulDivCtrl_isDiv;
  reg                 entries_0_uop_decoded_mulDivCtrl_isSigned;
  reg                 entries_0_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    entries_0_uop_decoded_memCtrl_size;
  reg                 entries_0_uop_decoded_memCtrl_isSignedLoad;
  reg                 entries_0_uop_decoded_memCtrl_isStore;
  reg                 entries_0_uop_decoded_memCtrl_isLoadLinked;
  reg                 entries_0_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    entries_0_uop_decoded_memCtrl_atomicOp;
  reg                 entries_0_uop_decoded_memCtrl_isFence;
  reg        [7:0]    entries_0_uop_decoded_memCtrl_fenceMode;
  reg                 entries_0_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    entries_0_uop_decoded_memCtrl_cacheOpType;
  reg                 entries_0_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    entries_0_uop_decoded_branchCtrl_condition;
  reg                 entries_0_uop_decoded_branchCtrl_isJump;
  reg                 entries_0_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    entries_0_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    entries_0_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 entries_0_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    entries_0_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    entries_0_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    entries_0_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    entries_0_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    entries_0_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    entries_0_uop_decoded_fpuCtrl_roundingMode;
  reg                 entries_0_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 entries_0_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 entries_0_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    entries_0_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   entries_0_uop_decoded_csrCtrl_csrAddr;
  reg                 entries_0_uop_decoded_csrCtrl_isWrite;
  reg                 entries_0_uop_decoded_csrCtrl_isRead;
  reg                 entries_0_uop_decoded_csrCtrl_isExchange;
  reg                 entries_0_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   entries_0_uop_decoded_sysCtrl_sysCode;
  reg                 entries_0_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 entries_0_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    entries_0_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    entries_0_uop_decoded_decodeExceptionCode;
  reg                 entries_0_uop_decoded_hasDecodeException;
  reg                 entries_0_uop_decoded_isMicrocode;
  reg        [7:0]    entries_0_uop_decoded_microcodeEntry;
  reg                 entries_0_uop_decoded_isSerializing;
  reg                 entries_0_uop_decoded_isBranchOrJump;
  reg                 entries_0_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   entries_0_uop_decoded_branchPrediction_target;
  reg                 entries_0_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    entries_0_uop_rename_physSrc1_idx;
  reg                 entries_0_uop_rename_physSrc1IsFpr;
  reg        [5:0]    entries_0_uop_rename_physSrc2_idx;
  reg                 entries_0_uop_rename_physSrc2IsFpr;
  reg        [5:0]    entries_0_uop_rename_physDest_idx;
  reg                 entries_0_uop_rename_physDestIsFpr;
  reg        [5:0]    entries_0_uop_rename_oldPhysDest_idx;
  reg                 entries_0_uop_rename_oldPhysDestIsFpr;
  reg                 entries_0_uop_rename_allocatesPhysDest;
  reg                 entries_0_uop_rename_writesToPhysReg;
  reg        [3:0]    entries_0_uop_robPtr;
  reg        [15:0]   entries_0_uop_uniqueId;
  reg                 entries_0_uop_dispatched;
  reg                 entries_0_uop_executed;
  reg                 entries_0_uop_hasException;
  reg        [7:0]    entries_0_uop_exceptionCode;
  reg        [3:0]    entries_0_robPtr;
  reg        [5:0]    entries_0_physDest_idx;
  reg                 entries_0_physDestIsFpr;
  reg                 entries_0_writesToPhysReg;
  reg                 entries_0_useSrc1;
  reg        [31:0]   entries_0_src1Data;
  reg        [5:0]    entries_0_src1Tag;
  reg                 entries_0_src1Ready;
  reg                 entries_0_src1IsFpr;
  reg                 entries_0_useSrc2;
  reg        [31:0]   entries_0_src2Data;
  reg        [5:0]    entries_0_src2Tag;
  reg                 entries_0_src2Ready;
  reg                 entries_0_src2IsFpr;
  reg                 entries_0_mulDivCtrl_valid;
  reg                 entries_0_mulDivCtrl_isDiv;
  reg                 entries_0_mulDivCtrl_isSigned;
  reg                 entries_0_mulDivCtrl_isWordOp;
  reg        [31:0]   entries_1_uop_decoded_pc;
  reg                 entries_1_uop_decoded_isValid;
  reg        [4:0]    entries_1_uop_decoded_uopCode;
  reg        [3:0]    entries_1_uop_decoded_exeUnit;
  reg        [1:0]    entries_1_uop_decoded_isa;
  reg        [4:0]    entries_1_uop_decoded_archDest_idx;
  reg        [1:0]    entries_1_uop_decoded_archDest_rtype;
  reg                 entries_1_uop_decoded_writeArchDestEn;
  reg        [4:0]    entries_1_uop_decoded_archSrc1_idx;
  reg        [1:0]    entries_1_uop_decoded_archSrc1_rtype;
  reg                 entries_1_uop_decoded_useArchSrc1;
  reg        [4:0]    entries_1_uop_decoded_archSrc2_idx;
  reg        [1:0]    entries_1_uop_decoded_archSrc2_rtype;
  reg                 entries_1_uop_decoded_useArchSrc2;
  reg                 entries_1_uop_decoded_usePcForAddr;
  reg        [31:0]   entries_1_uop_decoded_imm;
  reg        [2:0]    entries_1_uop_decoded_immUsage;
  reg                 entries_1_uop_decoded_aluCtrl_valid;
  reg                 entries_1_uop_decoded_aluCtrl_isSub;
  reg                 entries_1_uop_decoded_aluCtrl_isAdd;
  reg                 entries_1_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    entries_1_uop_decoded_aluCtrl_logicOp;
  reg                 entries_1_uop_decoded_shiftCtrl_valid;
  reg                 entries_1_uop_decoded_shiftCtrl_isRight;
  reg                 entries_1_uop_decoded_shiftCtrl_isArithmetic;
  reg                 entries_1_uop_decoded_shiftCtrl_isRotate;
  reg                 entries_1_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 entries_1_uop_decoded_mulDivCtrl_valid;
  reg                 entries_1_uop_decoded_mulDivCtrl_isDiv;
  reg                 entries_1_uop_decoded_mulDivCtrl_isSigned;
  reg                 entries_1_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    entries_1_uop_decoded_memCtrl_size;
  reg                 entries_1_uop_decoded_memCtrl_isSignedLoad;
  reg                 entries_1_uop_decoded_memCtrl_isStore;
  reg                 entries_1_uop_decoded_memCtrl_isLoadLinked;
  reg                 entries_1_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    entries_1_uop_decoded_memCtrl_atomicOp;
  reg                 entries_1_uop_decoded_memCtrl_isFence;
  reg        [7:0]    entries_1_uop_decoded_memCtrl_fenceMode;
  reg                 entries_1_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    entries_1_uop_decoded_memCtrl_cacheOpType;
  reg                 entries_1_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    entries_1_uop_decoded_branchCtrl_condition;
  reg                 entries_1_uop_decoded_branchCtrl_isJump;
  reg                 entries_1_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    entries_1_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    entries_1_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 entries_1_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    entries_1_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    entries_1_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    entries_1_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    entries_1_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    entries_1_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    entries_1_uop_decoded_fpuCtrl_roundingMode;
  reg                 entries_1_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 entries_1_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 entries_1_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    entries_1_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   entries_1_uop_decoded_csrCtrl_csrAddr;
  reg                 entries_1_uop_decoded_csrCtrl_isWrite;
  reg                 entries_1_uop_decoded_csrCtrl_isRead;
  reg                 entries_1_uop_decoded_csrCtrl_isExchange;
  reg                 entries_1_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   entries_1_uop_decoded_sysCtrl_sysCode;
  reg                 entries_1_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 entries_1_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    entries_1_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    entries_1_uop_decoded_decodeExceptionCode;
  reg                 entries_1_uop_decoded_hasDecodeException;
  reg                 entries_1_uop_decoded_isMicrocode;
  reg        [7:0]    entries_1_uop_decoded_microcodeEntry;
  reg                 entries_1_uop_decoded_isSerializing;
  reg                 entries_1_uop_decoded_isBranchOrJump;
  reg                 entries_1_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   entries_1_uop_decoded_branchPrediction_target;
  reg                 entries_1_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    entries_1_uop_rename_physSrc1_idx;
  reg                 entries_1_uop_rename_physSrc1IsFpr;
  reg        [5:0]    entries_1_uop_rename_physSrc2_idx;
  reg                 entries_1_uop_rename_physSrc2IsFpr;
  reg        [5:0]    entries_1_uop_rename_physDest_idx;
  reg                 entries_1_uop_rename_physDestIsFpr;
  reg        [5:0]    entries_1_uop_rename_oldPhysDest_idx;
  reg                 entries_1_uop_rename_oldPhysDestIsFpr;
  reg                 entries_1_uop_rename_allocatesPhysDest;
  reg                 entries_1_uop_rename_writesToPhysReg;
  reg        [3:0]    entries_1_uop_robPtr;
  reg        [15:0]   entries_1_uop_uniqueId;
  reg                 entries_1_uop_dispatched;
  reg                 entries_1_uop_executed;
  reg                 entries_1_uop_hasException;
  reg        [7:0]    entries_1_uop_exceptionCode;
  reg        [3:0]    entries_1_robPtr;
  reg        [5:0]    entries_1_physDest_idx;
  reg                 entries_1_physDestIsFpr;
  reg                 entries_1_writesToPhysReg;
  reg                 entries_1_useSrc1;
  reg        [31:0]   entries_1_src1Data;
  reg        [5:0]    entries_1_src1Tag;
  reg                 entries_1_src1Ready;
  reg                 entries_1_src1IsFpr;
  reg                 entries_1_useSrc2;
  reg        [31:0]   entries_1_src2Data;
  reg        [5:0]    entries_1_src2Tag;
  reg                 entries_1_src2Ready;
  reg                 entries_1_src2IsFpr;
  reg                 entries_1_mulDivCtrl_valid;
  reg                 entries_1_mulDivCtrl_isDiv;
  reg                 entries_1_mulDivCtrl_isSigned;
  reg                 entries_1_mulDivCtrl_isWordOp;
  reg        [31:0]   entries_2_uop_decoded_pc;
  reg                 entries_2_uop_decoded_isValid;
  reg        [4:0]    entries_2_uop_decoded_uopCode;
  reg        [3:0]    entries_2_uop_decoded_exeUnit;
  reg        [1:0]    entries_2_uop_decoded_isa;
  reg        [4:0]    entries_2_uop_decoded_archDest_idx;
  reg        [1:0]    entries_2_uop_decoded_archDest_rtype;
  reg                 entries_2_uop_decoded_writeArchDestEn;
  reg        [4:0]    entries_2_uop_decoded_archSrc1_idx;
  reg        [1:0]    entries_2_uop_decoded_archSrc1_rtype;
  reg                 entries_2_uop_decoded_useArchSrc1;
  reg        [4:0]    entries_2_uop_decoded_archSrc2_idx;
  reg        [1:0]    entries_2_uop_decoded_archSrc2_rtype;
  reg                 entries_2_uop_decoded_useArchSrc2;
  reg                 entries_2_uop_decoded_usePcForAddr;
  reg        [31:0]   entries_2_uop_decoded_imm;
  reg        [2:0]    entries_2_uop_decoded_immUsage;
  reg                 entries_2_uop_decoded_aluCtrl_valid;
  reg                 entries_2_uop_decoded_aluCtrl_isSub;
  reg                 entries_2_uop_decoded_aluCtrl_isAdd;
  reg                 entries_2_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    entries_2_uop_decoded_aluCtrl_logicOp;
  reg                 entries_2_uop_decoded_shiftCtrl_valid;
  reg                 entries_2_uop_decoded_shiftCtrl_isRight;
  reg                 entries_2_uop_decoded_shiftCtrl_isArithmetic;
  reg                 entries_2_uop_decoded_shiftCtrl_isRotate;
  reg                 entries_2_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 entries_2_uop_decoded_mulDivCtrl_valid;
  reg                 entries_2_uop_decoded_mulDivCtrl_isDiv;
  reg                 entries_2_uop_decoded_mulDivCtrl_isSigned;
  reg                 entries_2_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    entries_2_uop_decoded_memCtrl_size;
  reg                 entries_2_uop_decoded_memCtrl_isSignedLoad;
  reg                 entries_2_uop_decoded_memCtrl_isStore;
  reg                 entries_2_uop_decoded_memCtrl_isLoadLinked;
  reg                 entries_2_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    entries_2_uop_decoded_memCtrl_atomicOp;
  reg                 entries_2_uop_decoded_memCtrl_isFence;
  reg        [7:0]    entries_2_uop_decoded_memCtrl_fenceMode;
  reg                 entries_2_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    entries_2_uop_decoded_memCtrl_cacheOpType;
  reg                 entries_2_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    entries_2_uop_decoded_branchCtrl_condition;
  reg                 entries_2_uop_decoded_branchCtrl_isJump;
  reg                 entries_2_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    entries_2_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    entries_2_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 entries_2_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    entries_2_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    entries_2_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    entries_2_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    entries_2_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    entries_2_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    entries_2_uop_decoded_fpuCtrl_roundingMode;
  reg                 entries_2_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 entries_2_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 entries_2_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    entries_2_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   entries_2_uop_decoded_csrCtrl_csrAddr;
  reg                 entries_2_uop_decoded_csrCtrl_isWrite;
  reg                 entries_2_uop_decoded_csrCtrl_isRead;
  reg                 entries_2_uop_decoded_csrCtrl_isExchange;
  reg                 entries_2_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   entries_2_uop_decoded_sysCtrl_sysCode;
  reg                 entries_2_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 entries_2_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    entries_2_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    entries_2_uop_decoded_decodeExceptionCode;
  reg                 entries_2_uop_decoded_hasDecodeException;
  reg                 entries_2_uop_decoded_isMicrocode;
  reg        [7:0]    entries_2_uop_decoded_microcodeEntry;
  reg                 entries_2_uop_decoded_isSerializing;
  reg                 entries_2_uop_decoded_isBranchOrJump;
  reg                 entries_2_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   entries_2_uop_decoded_branchPrediction_target;
  reg                 entries_2_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    entries_2_uop_rename_physSrc1_idx;
  reg                 entries_2_uop_rename_physSrc1IsFpr;
  reg        [5:0]    entries_2_uop_rename_physSrc2_idx;
  reg                 entries_2_uop_rename_physSrc2IsFpr;
  reg        [5:0]    entries_2_uop_rename_physDest_idx;
  reg                 entries_2_uop_rename_physDestIsFpr;
  reg        [5:0]    entries_2_uop_rename_oldPhysDest_idx;
  reg                 entries_2_uop_rename_oldPhysDestIsFpr;
  reg                 entries_2_uop_rename_allocatesPhysDest;
  reg                 entries_2_uop_rename_writesToPhysReg;
  reg        [3:0]    entries_2_uop_robPtr;
  reg        [15:0]   entries_2_uop_uniqueId;
  reg                 entries_2_uop_dispatched;
  reg                 entries_2_uop_executed;
  reg                 entries_2_uop_hasException;
  reg        [7:0]    entries_2_uop_exceptionCode;
  reg        [3:0]    entries_2_robPtr;
  reg        [5:0]    entries_2_physDest_idx;
  reg                 entries_2_physDestIsFpr;
  reg                 entries_2_writesToPhysReg;
  reg                 entries_2_useSrc1;
  reg        [31:0]   entries_2_src1Data;
  reg        [5:0]    entries_2_src1Tag;
  reg                 entries_2_src1Ready;
  reg                 entries_2_src1IsFpr;
  reg                 entries_2_useSrc2;
  reg        [31:0]   entries_2_src2Data;
  reg        [5:0]    entries_2_src2Tag;
  reg                 entries_2_src2Ready;
  reg                 entries_2_src2IsFpr;
  reg                 entries_2_mulDivCtrl_valid;
  reg                 entries_2_mulDivCtrl_isDiv;
  reg                 entries_2_mulDivCtrl_isSigned;
  reg                 entries_2_mulDivCtrl_isWordOp;
  reg        [31:0]   entries_3_uop_decoded_pc;
  reg                 entries_3_uop_decoded_isValid;
  reg        [4:0]    entries_3_uop_decoded_uopCode;
  reg        [3:0]    entries_3_uop_decoded_exeUnit;
  reg        [1:0]    entries_3_uop_decoded_isa;
  reg        [4:0]    entries_3_uop_decoded_archDest_idx;
  reg        [1:0]    entries_3_uop_decoded_archDest_rtype;
  reg                 entries_3_uop_decoded_writeArchDestEn;
  reg        [4:0]    entries_3_uop_decoded_archSrc1_idx;
  reg        [1:0]    entries_3_uop_decoded_archSrc1_rtype;
  reg                 entries_3_uop_decoded_useArchSrc1;
  reg        [4:0]    entries_3_uop_decoded_archSrc2_idx;
  reg        [1:0]    entries_3_uop_decoded_archSrc2_rtype;
  reg                 entries_3_uop_decoded_useArchSrc2;
  reg                 entries_3_uop_decoded_usePcForAddr;
  reg        [31:0]   entries_3_uop_decoded_imm;
  reg        [2:0]    entries_3_uop_decoded_immUsage;
  reg                 entries_3_uop_decoded_aluCtrl_valid;
  reg                 entries_3_uop_decoded_aluCtrl_isSub;
  reg                 entries_3_uop_decoded_aluCtrl_isAdd;
  reg                 entries_3_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    entries_3_uop_decoded_aluCtrl_logicOp;
  reg                 entries_3_uop_decoded_shiftCtrl_valid;
  reg                 entries_3_uop_decoded_shiftCtrl_isRight;
  reg                 entries_3_uop_decoded_shiftCtrl_isArithmetic;
  reg                 entries_3_uop_decoded_shiftCtrl_isRotate;
  reg                 entries_3_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 entries_3_uop_decoded_mulDivCtrl_valid;
  reg                 entries_3_uop_decoded_mulDivCtrl_isDiv;
  reg                 entries_3_uop_decoded_mulDivCtrl_isSigned;
  reg                 entries_3_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    entries_3_uop_decoded_memCtrl_size;
  reg                 entries_3_uop_decoded_memCtrl_isSignedLoad;
  reg                 entries_3_uop_decoded_memCtrl_isStore;
  reg                 entries_3_uop_decoded_memCtrl_isLoadLinked;
  reg                 entries_3_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    entries_3_uop_decoded_memCtrl_atomicOp;
  reg                 entries_3_uop_decoded_memCtrl_isFence;
  reg        [7:0]    entries_3_uop_decoded_memCtrl_fenceMode;
  reg                 entries_3_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    entries_3_uop_decoded_memCtrl_cacheOpType;
  reg                 entries_3_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    entries_3_uop_decoded_branchCtrl_condition;
  reg                 entries_3_uop_decoded_branchCtrl_isJump;
  reg                 entries_3_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    entries_3_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    entries_3_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 entries_3_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    entries_3_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    entries_3_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    entries_3_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    entries_3_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    entries_3_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    entries_3_uop_decoded_fpuCtrl_roundingMode;
  reg                 entries_3_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 entries_3_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 entries_3_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    entries_3_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   entries_3_uop_decoded_csrCtrl_csrAddr;
  reg                 entries_3_uop_decoded_csrCtrl_isWrite;
  reg                 entries_3_uop_decoded_csrCtrl_isRead;
  reg                 entries_3_uop_decoded_csrCtrl_isExchange;
  reg                 entries_3_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   entries_3_uop_decoded_sysCtrl_sysCode;
  reg                 entries_3_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 entries_3_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    entries_3_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    entries_3_uop_decoded_decodeExceptionCode;
  reg                 entries_3_uop_decoded_hasDecodeException;
  reg                 entries_3_uop_decoded_isMicrocode;
  reg        [7:0]    entries_3_uop_decoded_microcodeEntry;
  reg                 entries_3_uop_decoded_isSerializing;
  reg                 entries_3_uop_decoded_isBranchOrJump;
  reg                 entries_3_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   entries_3_uop_decoded_branchPrediction_target;
  reg                 entries_3_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    entries_3_uop_rename_physSrc1_idx;
  reg                 entries_3_uop_rename_physSrc1IsFpr;
  reg        [5:0]    entries_3_uop_rename_physSrc2_idx;
  reg                 entries_3_uop_rename_physSrc2IsFpr;
  reg        [5:0]    entries_3_uop_rename_physDest_idx;
  reg                 entries_3_uop_rename_physDestIsFpr;
  reg        [5:0]    entries_3_uop_rename_oldPhysDest_idx;
  reg                 entries_3_uop_rename_oldPhysDestIsFpr;
  reg                 entries_3_uop_rename_allocatesPhysDest;
  reg                 entries_3_uop_rename_writesToPhysReg;
  reg        [3:0]    entries_3_uop_robPtr;
  reg        [15:0]   entries_3_uop_uniqueId;
  reg                 entries_3_uop_dispatched;
  reg                 entries_3_uop_executed;
  reg                 entries_3_uop_hasException;
  reg        [7:0]    entries_3_uop_exceptionCode;
  reg        [3:0]    entries_3_robPtr;
  reg        [5:0]    entries_3_physDest_idx;
  reg                 entries_3_physDestIsFpr;
  reg                 entries_3_writesToPhysReg;
  reg                 entries_3_useSrc1;
  reg        [31:0]   entries_3_src1Data;
  reg        [5:0]    entries_3_src1Tag;
  reg                 entries_3_src1Ready;
  reg                 entries_3_src1IsFpr;
  reg                 entries_3_useSrc2;
  reg        [31:0]   entries_3_src2Data;
  reg        [5:0]    entries_3_src2Tag;
  reg                 entries_3_src2Ready;
  reg                 entries_3_src2IsFpr;
  reg                 entries_3_mulDivCtrl_valid;
  reg                 entries_3_mulDivCtrl_isDiv;
  reg                 entries_3_mulDivCtrl_isSigned;
  reg                 entries_3_mulDivCtrl_isWordOp;
  reg                 entryValids_0;
  reg                 entryValids_1;
  reg                 entryValids_2;
  reg                 entryValids_3;
  wire                io_issueOut_fire;
  wire                localWakeupValid;
  reg        [3:0]    wokeUpSrc1Mask;
  reg        [3:0]    wokeUpSrc2Mask;
  wire                _zz_when_IssueQueueComponent_l103;
  wire                _zz_when_IssueQueueComponent_l106;
  wire                when_IssueQueueComponent_l103;
  wire                when_IssueQueueComponent_l106;
  wire                when_IssueQueueComponent_l113;
  wire                when_IssueQueueComponent_l116;
  wire                when_IssueQueueComponent_l113_1;
  wire                when_IssueQueueComponent_l116_1;
  wire                when_IssueQueueComponent_l113_2;
  wire                when_IssueQueueComponent_l116_2;
  wire                when_IssueQueueComponent_l113_3;
  wire                when_IssueQueueComponent_l116_3;
  wire                when_IssueQueueComponent_l113_4;
  wire                when_IssueQueueComponent_l116_4;
  wire                _zz_when_IssueQueueComponent_l103_1;
  wire                _zz_when_IssueQueueComponent_l106_1;
  wire                when_IssueQueueComponent_l103_1;
  wire                when_IssueQueueComponent_l106_1;
  wire                when_IssueQueueComponent_l113_5;
  wire                when_IssueQueueComponent_l116_5;
  wire                when_IssueQueueComponent_l113_6;
  wire                when_IssueQueueComponent_l116_6;
  wire                when_IssueQueueComponent_l113_7;
  wire                when_IssueQueueComponent_l116_7;
  wire                when_IssueQueueComponent_l113_8;
  wire                when_IssueQueueComponent_l116_8;
  wire                when_IssueQueueComponent_l113_9;
  wire                when_IssueQueueComponent_l116_9;
  wire                _zz_when_IssueQueueComponent_l103_2;
  wire                _zz_when_IssueQueueComponent_l106_2;
  wire                when_IssueQueueComponent_l103_2;
  wire                when_IssueQueueComponent_l106_2;
  wire                when_IssueQueueComponent_l113_10;
  wire                when_IssueQueueComponent_l116_10;
  wire                when_IssueQueueComponent_l113_11;
  wire                when_IssueQueueComponent_l116_11;
  wire                when_IssueQueueComponent_l113_12;
  wire                when_IssueQueueComponent_l116_12;
  wire                when_IssueQueueComponent_l113_13;
  wire                when_IssueQueueComponent_l116_13;
  wire                when_IssueQueueComponent_l113_14;
  wire                when_IssueQueueComponent_l116_14;
  wire                _zz_when_IssueQueueComponent_l103_3;
  wire                _zz_when_IssueQueueComponent_l106_3;
  wire                when_IssueQueueComponent_l103_3;
  wire                when_IssueQueueComponent_l106_3;
  wire                when_IssueQueueComponent_l113_15;
  wire                when_IssueQueueComponent_l116_15;
  wire                when_IssueQueueComponent_l113_16;
  wire                when_IssueQueueComponent_l116_16;
  wire                when_IssueQueueComponent_l113_17;
  wire                when_IssueQueueComponent_l116_17;
  wire                when_IssueQueueComponent_l113_18;
  wire                when_IssueQueueComponent_l116_18;
  wire                when_IssueQueueComponent_l113_19;
  wire                when_IssueQueueComponent_l116_19;
  wire                entriesReadyToIssue_0;
  wire                entriesReadyToIssue_1;
  wire                entriesReadyToIssue_2;
  wire                entriesReadyToIssue_3;
  wire       [3:0]    issueRequestMask;
  wire       [3:0]    issueRequestMask_ohFirst_input;
  wire       [3:0]    issueRequestMask_ohFirst_masked;
  wire       [3:0]    issueRequestOh;
  wire                _zz_issueIdx;
  wire                _zz_issueIdx_1;
  wire                _zz_issueIdx_2;
  wire       [1:0]    issueIdx;
  wire       [4:0]    _zz_io_issueOut_payload_uop_decoded_uopCode;
  wire       [3:0]    _zz_io_issueOut_payload_uop_decoded_exeUnit;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_isa;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_archDest_rtype;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype;
  wire       [2:0]    _zz_io_issueOut_payload_uop_decoded_immUsage;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_memCtrl_size;
  wire       [4:0]    _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest;
  wire       [1:0]    _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode;
  wire       [3:0]    freeSlotsMask;
  wire                hasSpaceForNewEntry;
  reg        [3:0]    firedSlotMask;
  wire       [3:0]    _zz_allocationMask;
  wire       [3:0]    allocationMask;
  wire                _zz_allocateIdx;
  wire                _zz_allocateIdx_1;
  wire                _zz_allocateIdx_2;
  wire       [1:0]    allocateIdx;
  reg        [31:0]   entriesNext_0_uop_decoded_pc;
  reg                 entriesNext_0_uop_decoded_isValid;
  reg        [4:0]    entriesNext_0_uop_decoded_uopCode;
  reg        [3:0]    entriesNext_0_uop_decoded_exeUnit;
  reg        [1:0]    entriesNext_0_uop_decoded_isa;
  reg        [4:0]    entriesNext_0_uop_decoded_archDest_idx;
  reg        [1:0]    entriesNext_0_uop_decoded_archDest_rtype;
  reg                 entriesNext_0_uop_decoded_writeArchDestEn;
  reg        [4:0]    entriesNext_0_uop_decoded_archSrc1_idx;
  reg        [1:0]    entriesNext_0_uop_decoded_archSrc1_rtype;
  reg                 entriesNext_0_uop_decoded_useArchSrc1;
  reg        [4:0]    entriesNext_0_uop_decoded_archSrc2_idx;
  reg        [1:0]    entriesNext_0_uop_decoded_archSrc2_rtype;
  reg                 entriesNext_0_uop_decoded_useArchSrc2;
  reg                 entriesNext_0_uop_decoded_usePcForAddr;
  reg        [31:0]   entriesNext_0_uop_decoded_imm;
  reg        [2:0]    entriesNext_0_uop_decoded_immUsage;
  reg                 entriesNext_0_uop_decoded_aluCtrl_valid;
  reg                 entriesNext_0_uop_decoded_aluCtrl_isSub;
  reg                 entriesNext_0_uop_decoded_aluCtrl_isAdd;
  reg                 entriesNext_0_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    entriesNext_0_uop_decoded_aluCtrl_logicOp;
  reg                 entriesNext_0_uop_decoded_shiftCtrl_valid;
  reg                 entriesNext_0_uop_decoded_shiftCtrl_isRight;
  reg                 entriesNext_0_uop_decoded_shiftCtrl_isArithmetic;
  reg                 entriesNext_0_uop_decoded_shiftCtrl_isRotate;
  reg                 entriesNext_0_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 entriesNext_0_uop_decoded_mulDivCtrl_valid;
  reg                 entriesNext_0_uop_decoded_mulDivCtrl_isDiv;
  reg                 entriesNext_0_uop_decoded_mulDivCtrl_isSigned;
  reg                 entriesNext_0_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    entriesNext_0_uop_decoded_memCtrl_size;
  reg                 entriesNext_0_uop_decoded_memCtrl_isSignedLoad;
  reg                 entriesNext_0_uop_decoded_memCtrl_isStore;
  reg                 entriesNext_0_uop_decoded_memCtrl_isLoadLinked;
  reg                 entriesNext_0_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    entriesNext_0_uop_decoded_memCtrl_atomicOp;
  reg                 entriesNext_0_uop_decoded_memCtrl_isFence;
  reg        [7:0]    entriesNext_0_uop_decoded_memCtrl_fenceMode;
  reg                 entriesNext_0_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    entriesNext_0_uop_decoded_memCtrl_cacheOpType;
  reg                 entriesNext_0_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    entriesNext_0_uop_decoded_branchCtrl_condition;
  reg                 entriesNext_0_uop_decoded_branchCtrl_isJump;
  reg                 entriesNext_0_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    entriesNext_0_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 entriesNext_0_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    entriesNext_0_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    entriesNext_0_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    entriesNext_0_uop_decoded_fpuCtrl_roundingMode;
  reg                 entriesNext_0_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 entriesNext_0_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 entriesNext_0_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    entriesNext_0_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   entriesNext_0_uop_decoded_csrCtrl_csrAddr;
  reg                 entriesNext_0_uop_decoded_csrCtrl_isWrite;
  reg                 entriesNext_0_uop_decoded_csrCtrl_isRead;
  reg                 entriesNext_0_uop_decoded_csrCtrl_isExchange;
  reg                 entriesNext_0_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   entriesNext_0_uop_decoded_sysCtrl_sysCode;
  reg                 entriesNext_0_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 entriesNext_0_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    entriesNext_0_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    entriesNext_0_uop_decoded_decodeExceptionCode;
  reg                 entriesNext_0_uop_decoded_hasDecodeException;
  reg                 entriesNext_0_uop_decoded_isMicrocode;
  reg        [7:0]    entriesNext_0_uop_decoded_microcodeEntry;
  reg                 entriesNext_0_uop_decoded_isSerializing;
  reg                 entriesNext_0_uop_decoded_isBranchOrJump;
  reg                 entriesNext_0_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   entriesNext_0_uop_decoded_branchPrediction_target;
  reg                 entriesNext_0_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    entriesNext_0_uop_rename_physSrc1_idx;
  reg                 entriesNext_0_uop_rename_physSrc1IsFpr;
  reg        [5:0]    entriesNext_0_uop_rename_physSrc2_idx;
  reg                 entriesNext_0_uop_rename_physSrc2IsFpr;
  reg        [5:0]    entriesNext_0_uop_rename_physDest_idx;
  reg                 entriesNext_0_uop_rename_physDestIsFpr;
  reg        [5:0]    entriesNext_0_uop_rename_oldPhysDest_idx;
  reg                 entriesNext_0_uop_rename_oldPhysDestIsFpr;
  reg                 entriesNext_0_uop_rename_allocatesPhysDest;
  reg                 entriesNext_0_uop_rename_writesToPhysReg;
  reg        [3:0]    entriesNext_0_uop_robPtr;
  reg        [15:0]   entriesNext_0_uop_uniqueId;
  reg                 entriesNext_0_uop_dispatched;
  reg                 entriesNext_0_uop_executed;
  reg                 entriesNext_0_uop_hasException;
  reg        [7:0]    entriesNext_0_uop_exceptionCode;
  reg        [3:0]    entriesNext_0_robPtr;
  reg        [5:0]    entriesNext_0_physDest_idx;
  reg                 entriesNext_0_physDestIsFpr;
  reg                 entriesNext_0_writesToPhysReg;
  reg                 entriesNext_0_useSrc1;
  reg        [31:0]   entriesNext_0_src1Data;
  reg        [5:0]    entriesNext_0_src1Tag;
  reg                 entriesNext_0_src1Ready;
  reg                 entriesNext_0_src1IsFpr;
  reg                 entriesNext_0_useSrc2;
  reg        [31:0]   entriesNext_0_src2Data;
  reg        [5:0]    entriesNext_0_src2Tag;
  reg                 entriesNext_0_src2Ready;
  reg                 entriesNext_0_src2IsFpr;
  reg                 entriesNext_0_mulDivCtrl_valid;
  reg                 entriesNext_0_mulDivCtrl_isDiv;
  reg                 entriesNext_0_mulDivCtrl_isSigned;
  reg                 entriesNext_0_mulDivCtrl_isWordOp;
  reg        [31:0]   entriesNext_1_uop_decoded_pc;
  reg                 entriesNext_1_uop_decoded_isValid;
  reg        [4:0]    entriesNext_1_uop_decoded_uopCode;
  reg        [3:0]    entriesNext_1_uop_decoded_exeUnit;
  reg        [1:0]    entriesNext_1_uop_decoded_isa;
  reg        [4:0]    entriesNext_1_uop_decoded_archDest_idx;
  reg        [1:0]    entriesNext_1_uop_decoded_archDest_rtype;
  reg                 entriesNext_1_uop_decoded_writeArchDestEn;
  reg        [4:0]    entriesNext_1_uop_decoded_archSrc1_idx;
  reg        [1:0]    entriesNext_1_uop_decoded_archSrc1_rtype;
  reg                 entriesNext_1_uop_decoded_useArchSrc1;
  reg        [4:0]    entriesNext_1_uop_decoded_archSrc2_idx;
  reg        [1:0]    entriesNext_1_uop_decoded_archSrc2_rtype;
  reg                 entriesNext_1_uop_decoded_useArchSrc2;
  reg                 entriesNext_1_uop_decoded_usePcForAddr;
  reg        [31:0]   entriesNext_1_uop_decoded_imm;
  reg        [2:0]    entriesNext_1_uop_decoded_immUsage;
  reg                 entriesNext_1_uop_decoded_aluCtrl_valid;
  reg                 entriesNext_1_uop_decoded_aluCtrl_isSub;
  reg                 entriesNext_1_uop_decoded_aluCtrl_isAdd;
  reg                 entriesNext_1_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    entriesNext_1_uop_decoded_aluCtrl_logicOp;
  reg                 entriesNext_1_uop_decoded_shiftCtrl_valid;
  reg                 entriesNext_1_uop_decoded_shiftCtrl_isRight;
  reg                 entriesNext_1_uop_decoded_shiftCtrl_isArithmetic;
  reg                 entriesNext_1_uop_decoded_shiftCtrl_isRotate;
  reg                 entriesNext_1_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 entriesNext_1_uop_decoded_mulDivCtrl_valid;
  reg                 entriesNext_1_uop_decoded_mulDivCtrl_isDiv;
  reg                 entriesNext_1_uop_decoded_mulDivCtrl_isSigned;
  reg                 entriesNext_1_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    entriesNext_1_uop_decoded_memCtrl_size;
  reg                 entriesNext_1_uop_decoded_memCtrl_isSignedLoad;
  reg                 entriesNext_1_uop_decoded_memCtrl_isStore;
  reg                 entriesNext_1_uop_decoded_memCtrl_isLoadLinked;
  reg                 entriesNext_1_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    entriesNext_1_uop_decoded_memCtrl_atomicOp;
  reg                 entriesNext_1_uop_decoded_memCtrl_isFence;
  reg        [7:0]    entriesNext_1_uop_decoded_memCtrl_fenceMode;
  reg                 entriesNext_1_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    entriesNext_1_uop_decoded_memCtrl_cacheOpType;
  reg                 entriesNext_1_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    entriesNext_1_uop_decoded_branchCtrl_condition;
  reg                 entriesNext_1_uop_decoded_branchCtrl_isJump;
  reg                 entriesNext_1_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    entriesNext_1_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 entriesNext_1_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    entriesNext_1_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    entriesNext_1_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    entriesNext_1_uop_decoded_fpuCtrl_roundingMode;
  reg                 entriesNext_1_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 entriesNext_1_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 entriesNext_1_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    entriesNext_1_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   entriesNext_1_uop_decoded_csrCtrl_csrAddr;
  reg                 entriesNext_1_uop_decoded_csrCtrl_isWrite;
  reg                 entriesNext_1_uop_decoded_csrCtrl_isRead;
  reg                 entriesNext_1_uop_decoded_csrCtrl_isExchange;
  reg                 entriesNext_1_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   entriesNext_1_uop_decoded_sysCtrl_sysCode;
  reg                 entriesNext_1_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 entriesNext_1_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    entriesNext_1_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    entriesNext_1_uop_decoded_decodeExceptionCode;
  reg                 entriesNext_1_uop_decoded_hasDecodeException;
  reg                 entriesNext_1_uop_decoded_isMicrocode;
  reg        [7:0]    entriesNext_1_uop_decoded_microcodeEntry;
  reg                 entriesNext_1_uop_decoded_isSerializing;
  reg                 entriesNext_1_uop_decoded_isBranchOrJump;
  reg                 entriesNext_1_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   entriesNext_1_uop_decoded_branchPrediction_target;
  reg                 entriesNext_1_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    entriesNext_1_uop_rename_physSrc1_idx;
  reg                 entriesNext_1_uop_rename_physSrc1IsFpr;
  reg        [5:0]    entriesNext_1_uop_rename_physSrc2_idx;
  reg                 entriesNext_1_uop_rename_physSrc2IsFpr;
  reg        [5:0]    entriesNext_1_uop_rename_physDest_idx;
  reg                 entriesNext_1_uop_rename_physDestIsFpr;
  reg        [5:0]    entriesNext_1_uop_rename_oldPhysDest_idx;
  reg                 entriesNext_1_uop_rename_oldPhysDestIsFpr;
  reg                 entriesNext_1_uop_rename_allocatesPhysDest;
  reg                 entriesNext_1_uop_rename_writesToPhysReg;
  reg        [3:0]    entriesNext_1_uop_robPtr;
  reg        [15:0]   entriesNext_1_uop_uniqueId;
  reg                 entriesNext_1_uop_dispatched;
  reg                 entriesNext_1_uop_executed;
  reg                 entriesNext_1_uop_hasException;
  reg        [7:0]    entriesNext_1_uop_exceptionCode;
  reg        [3:0]    entriesNext_1_robPtr;
  reg        [5:0]    entriesNext_1_physDest_idx;
  reg                 entriesNext_1_physDestIsFpr;
  reg                 entriesNext_1_writesToPhysReg;
  reg                 entriesNext_1_useSrc1;
  reg        [31:0]   entriesNext_1_src1Data;
  reg        [5:0]    entriesNext_1_src1Tag;
  reg                 entriesNext_1_src1Ready;
  reg                 entriesNext_1_src1IsFpr;
  reg                 entriesNext_1_useSrc2;
  reg        [31:0]   entriesNext_1_src2Data;
  reg        [5:0]    entriesNext_1_src2Tag;
  reg                 entriesNext_1_src2Ready;
  reg                 entriesNext_1_src2IsFpr;
  reg                 entriesNext_1_mulDivCtrl_valid;
  reg                 entriesNext_1_mulDivCtrl_isDiv;
  reg                 entriesNext_1_mulDivCtrl_isSigned;
  reg                 entriesNext_1_mulDivCtrl_isWordOp;
  reg        [31:0]   entriesNext_2_uop_decoded_pc;
  reg                 entriesNext_2_uop_decoded_isValid;
  reg        [4:0]    entriesNext_2_uop_decoded_uopCode;
  reg        [3:0]    entriesNext_2_uop_decoded_exeUnit;
  reg        [1:0]    entriesNext_2_uop_decoded_isa;
  reg        [4:0]    entriesNext_2_uop_decoded_archDest_idx;
  reg        [1:0]    entriesNext_2_uop_decoded_archDest_rtype;
  reg                 entriesNext_2_uop_decoded_writeArchDestEn;
  reg        [4:0]    entriesNext_2_uop_decoded_archSrc1_idx;
  reg        [1:0]    entriesNext_2_uop_decoded_archSrc1_rtype;
  reg                 entriesNext_2_uop_decoded_useArchSrc1;
  reg        [4:0]    entriesNext_2_uop_decoded_archSrc2_idx;
  reg        [1:0]    entriesNext_2_uop_decoded_archSrc2_rtype;
  reg                 entriesNext_2_uop_decoded_useArchSrc2;
  reg                 entriesNext_2_uop_decoded_usePcForAddr;
  reg        [31:0]   entriesNext_2_uop_decoded_imm;
  reg        [2:0]    entriesNext_2_uop_decoded_immUsage;
  reg                 entriesNext_2_uop_decoded_aluCtrl_valid;
  reg                 entriesNext_2_uop_decoded_aluCtrl_isSub;
  reg                 entriesNext_2_uop_decoded_aluCtrl_isAdd;
  reg                 entriesNext_2_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    entriesNext_2_uop_decoded_aluCtrl_logicOp;
  reg                 entriesNext_2_uop_decoded_shiftCtrl_valid;
  reg                 entriesNext_2_uop_decoded_shiftCtrl_isRight;
  reg                 entriesNext_2_uop_decoded_shiftCtrl_isArithmetic;
  reg                 entriesNext_2_uop_decoded_shiftCtrl_isRotate;
  reg                 entriesNext_2_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 entriesNext_2_uop_decoded_mulDivCtrl_valid;
  reg                 entriesNext_2_uop_decoded_mulDivCtrl_isDiv;
  reg                 entriesNext_2_uop_decoded_mulDivCtrl_isSigned;
  reg                 entriesNext_2_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    entriesNext_2_uop_decoded_memCtrl_size;
  reg                 entriesNext_2_uop_decoded_memCtrl_isSignedLoad;
  reg                 entriesNext_2_uop_decoded_memCtrl_isStore;
  reg                 entriesNext_2_uop_decoded_memCtrl_isLoadLinked;
  reg                 entriesNext_2_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    entriesNext_2_uop_decoded_memCtrl_atomicOp;
  reg                 entriesNext_2_uop_decoded_memCtrl_isFence;
  reg        [7:0]    entriesNext_2_uop_decoded_memCtrl_fenceMode;
  reg                 entriesNext_2_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    entriesNext_2_uop_decoded_memCtrl_cacheOpType;
  reg                 entriesNext_2_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    entriesNext_2_uop_decoded_branchCtrl_condition;
  reg                 entriesNext_2_uop_decoded_branchCtrl_isJump;
  reg                 entriesNext_2_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    entriesNext_2_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 entriesNext_2_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    entriesNext_2_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    entriesNext_2_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    entriesNext_2_uop_decoded_fpuCtrl_roundingMode;
  reg                 entriesNext_2_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 entriesNext_2_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 entriesNext_2_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    entriesNext_2_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   entriesNext_2_uop_decoded_csrCtrl_csrAddr;
  reg                 entriesNext_2_uop_decoded_csrCtrl_isWrite;
  reg                 entriesNext_2_uop_decoded_csrCtrl_isRead;
  reg                 entriesNext_2_uop_decoded_csrCtrl_isExchange;
  reg                 entriesNext_2_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   entriesNext_2_uop_decoded_sysCtrl_sysCode;
  reg                 entriesNext_2_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 entriesNext_2_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    entriesNext_2_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    entriesNext_2_uop_decoded_decodeExceptionCode;
  reg                 entriesNext_2_uop_decoded_hasDecodeException;
  reg                 entriesNext_2_uop_decoded_isMicrocode;
  reg        [7:0]    entriesNext_2_uop_decoded_microcodeEntry;
  reg                 entriesNext_2_uop_decoded_isSerializing;
  reg                 entriesNext_2_uop_decoded_isBranchOrJump;
  reg                 entriesNext_2_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   entriesNext_2_uop_decoded_branchPrediction_target;
  reg                 entriesNext_2_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    entriesNext_2_uop_rename_physSrc1_idx;
  reg                 entriesNext_2_uop_rename_physSrc1IsFpr;
  reg        [5:0]    entriesNext_2_uop_rename_physSrc2_idx;
  reg                 entriesNext_2_uop_rename_physSrc2IsFpr;
  reg        [5:0]    entriesNext_2_uop_rename_physDest_idx;
  reg                 entriesNext_2_uop_rename_physDestIsFpr;
  reg        [5:0]    entriesNext_2_uop_rename_oldPhysDest_idx;
  reg                 entriesNext_2_uop_rename_oldPhysDestIsFpr;
  reg                 entriesNext_2_uop_rename_allocatesPhysDest;
  reg                 entriesNext_2_uop_rename_writesToPhysReg;
  reg        [3:0]    entriesNext_2_uop_robPtr;
  reg        [15:0]   entriesNext_2_uop_uniqueId;
  reg                 entriesNext_2_uop_dispatched;
  reg                 entriesNext_2_uop_executed;
  reg                 entriesNext_2_uop_hasException;
  reg        [7:0]    entriesNext_2_uop_exceptionCode;
  reg        [3:0]    entriesNext_2_robPtr;
  reg        [5:0]    entriesNext_2_physDest_idx;
  reg                 entriesNext_2_physDestIsFpr;
  reg                 entriesNext_2_writesToPhysReg;
  reg                 entriesNext_2_useSrc1;
  reg        [31:0]   entriesNext_2_src1Data;
  reg        [5:0]    entriesNext_2_src1Tag;
  reg                 entriesNext_2_src1Ready;
  reg                 entriesNext_2_src1IsFpr;
  reg                 entriesNext_2_useSrc2;
  reg        [31:0]   entriesNext_2_src2Data;
  reg        [5:0]    entriesNext_2_src2Tag;
  reg                 entriesNext_2_src2Ready;
  reg                 entriesNext_2_src2IsFpr;
  reg                 entriesNext_2_mulDivCtrl_valid;
  reg                 entriesNext_2_mulDivCtrl_isDiv;
  reg                 entriesNext_2_mulDivCtrl_isSigned;
  reg                 entriesNext_2_mulDivCtrl_isWordOp;
  reg        [31:0]   entriesNext_3_uop_decoded_pc;
  reg                 entriesNext_3_uop_decoded_isValid;
  reg        [4:0]    entriesNext_3_uop_decoded_uopCode;
  reg        [3:0]    entriesNext_3_uop_decoded_exeUnit;
  reg        [1:0]    entriesNext_3_uop_decoded_isa;
  reg        [4:0]    entriesNext_3_uop_decoded_archDest_idx;
  reg        [1:0]    entriesNext_3_uop_decoded_archDest_rtype;
  reg                 entriesNext_3_uop_decoded_writeArchDestEn;
  reg        [4:0]    entriesNext_3_uop_decoded_archSrc1_idx;
  reg        [1:0]    entriesNext_3_uop_decoded_archSrc1_rtype;
  reg                 entriesNext_3_uop_decoded_useArchSrc1;
  reg        [4:0]    entriesNext_3_uop_decoded_archSrc2_idx;
  reg        [1:0]    entriesNext_3_uop_decoded_archSrc2_rtype;
  reg                 entriesNext_3_uop_decoded_useArchSrc2;
  reg                 entriesNext_3_uop_decoded_usePcForAddr;
  reg        [31:0]   entriesNext_3_uop_decoded_imm;
  reg        [2:0]    entriesNext_3_uop_decoded_immUsage;
  reg                 entriesNext_3_uop_decoded_aluCtrl_valid;
  reg                 entriesNext_3_uop_decoded_aluCtrl_isSub;
  reg                 entriesNext_3_uop_decoded_aluCtrl_isAdd;
  reg                 entriesNext_3_uop_decoded_aluCtrl_isSigned;
  reg        [1:0]    entriesNext_3_uop_decoded_aluCtrl_logicOp;
  reg                 entriesNext_3_uop_decoded_shiftCtrl_valid;
  reg                 entriesNext_3_uop_decoded_shiftCtrl_isRight;
  reg                 entriesNext_3_uop_decoded_shiftCtrl_isArithmetic;
  reg                 entriesNext_3_uop_decoded_shiftCtrl_isRotate;
  reg                 entriesNext_3_uop_decoded_shiftCtrl_isDoubleWord;
  reg                 entriesNext_3_uop_decoded_mulDivCtrl_valid;
  reg                 entriesNext_3_uop_decoded_mulDivCtrl_isDiv;
  reg                 entriesNext_3_uop_decoded_mulDivCtrl_isSigned;
  reg                 entriesNext_3_uop_decoded_mulDivCtrl_isWordOp;
  reg        [1:0]    entriesNext_3_uop_decoded_memCtrl_size;
  reg                 entriesNext_3_uop_decoded_memCtrl_isSignedLoad;
  reg                 entriesNext_3_uop_decoded_memCtrl_isStore;
  reg                 entriesNext_3_uop_decoded_memCtrl_isLoadLinked;
  reg                 entriesNext_3_uop_decoded_memCtrl_isStoreCond;
  reg        [4:0]    entriesNext_3_uop_decoded_memCtrl_atomicOp;
  reg                 entriesNext_3_uop_decoded_memCtrl_isFence;
  reg        [7:0]    entriesNext_3_uop_decoded_memCtrl_fenceMode;
  reg                 entriesNext_3_uop_decoded_memCtrl_isCacheOp;
  reg        [4:0]    entriesNext_3_uop_decoded_memCtrl_cacheOpType;
  reg                 entriesNext_3_uop_decoded_memCtrl_isPrefetch;
  reg        [4:0]    entriesNext_3_uop_decoded_branchCtrl_condition;
  reg                 entriesNext_3_uop_decoded_branchCtrl_isJump;
  reg                 entriesNext_3_uop_decoded_branchCtrl_isLink;
  reg        [4:0]    entriesNext_3_uop_decoded_branchCtrl_linkReg_idx;
  reg        [1:0]    entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype;
  reg                 entriesNext_3_uop_decoded_branchCtrl_isIndirect;
  reg        [2:0]    entriesNext_3_uop_decoded_branchCtrl_laCfIdx;
  reg        [3:0]    entriesNext_3_uop_decoded_fpuCtrl_opType;
  reg        [1:0]    entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1;
  reg        [1:0]    entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2;
  reg        [1:0]    entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest;
  reg        [2:0]    entriesNext_3_uop_decoded_fpuCtrl_roundingMode;
  reg                 entriesNext_3_uop_decoded_fpuCtrl_isIntegerDest;
  reg                 entriesNext_3_uop_decoded_fpuCtrl_isSignedCvt;
  reg                 entriesNext_3_uop_decoded_fpuCtrl_fmaNegSrc1;
  reg        [4:0]    entriesNext_3_uop_decoded_fpuCtrl_fcmpCond;
  reg        [13:0]   entriesNext_3_uop_decoded_csrCtrl_csrAddr;
  reg                 entriesNext_3_uop_decoded_csrCtrl_isWrite;
  reg                 entriesNext_3_uop_decoded_csrCtrl_isRead;
  reg                 entriesNext_3_uop_decoded_csrCtrl_isExchange;
  reg                 entriesNext_3_uop_decoded_csrCtrl_useUimmAsSrc;
  reg        [19:0]   entriesNext_3_uop_decoded_sysCtrl_sysCode;
  reg                 entriesNext_3_uop_decoded_sysCtrl_isExceptionReturn;
  reg                 entriesNext_3_uop_decoded_sysCtrl_isTlbOp;
  reg        [3:0]    entriesNext_3_uop_decoded_sysCtrl_tlbOpType;
  reg        [1:0]    entriesNext_3_uop_decoded_decodeExceptionCode;
  reg                 entriesNext_3_uop_decoded_hasDecodeException;
  reg                 entriesNext_3_uop_decoded_isMicrocode;
  reg        [7:0]    entriesNext_3_uop_decoded_microcodeEntry;
  reg                 entriesNext_3_uop_decoded_isSerializing;
  reg                 entriesNext_3_uop_decoded_isBranchOrJump;
  reg                 entriesNext_3_uop_decoded_branchPrediction_isTaken;
  reg        [31:0]   entriesNext_3_uop_decoded_branchPrediction_target;
  reg                 entriesNext_3_uop_decoded_branchPrediction_wasPredicted;
  reg        [5:0]    entriesNext_3_uop_rename_physSrc1_idx;
  reg                 entriesNext_3_uop_rename_physSrc1IsFpr;
  reg        [5:0]    entriesNext_3_uop_rename_physSrc2_idx;
  reg                 entriesNext_3_uop_rename_physSrc2IsFpr;
  reg        [5:0]    entriesNext_3_uop_rename_physDest_idx;
  reg                 entriesNext_3_uop_rename_physDestIsFpr;
  reg        [5:0]    entriesNext_3_uop_rename_oldPhysDest_idx;
  reg                 entriesNext_3_uop_rename_oldPhysDestIsFpr;
  reg                 entriesNext_3_uop_rename_allocatesPhysDest;
  reg                 entriesNext_3_uop_rename_writesToPhysReg;
  reg        [3:0]    entriesNext_3_uop_robPtr;
  reg        [15:0]   entriesNext_3_uop_uniqueId;
  reg                 entriesNext_3_uop_dispatched;
  reg                 entriesNext_3_uop_executed;
  reg                 entriesNext_3_uop_hasException;
  reg        [7:0]    entriesNext_3_uop_exceptionCode;
  reg        [3:0]    entriesNext_3_robPtr;
  reg        [5:0]    entriesNext_3_physDest_idx;
  reg                 entriesNext_3_physDestIsFpr;
  reg                 entriesNext_3_writesToPhysReg;
  reg                 entriesNext_3_useSrc1;
  reg        [31:0]   entriesNext_3_src1Data;
  reg        [5:0]    entriesNext_3_src1Tag;
  reg                 entriesNext_3_src1Ready;
  reg                 entriesNext_3_src1IsFpr;
  reg                 entriesNext_3_useSrc2;
  reg        [31:0]   entriesNext_3_src2Data;
  reg        [5:0]    entriesNext_3_src2Tag;
  reg                 entriesNext_3_src2Ready;
  reg                 entriesNext_3_src2IsFpr;
  reg                 entriesNext_3_mulDivCtrl_valid;
  reg                 entriesNext_3_mulDivCtrl_isDiv;
  reg                 entriesNext_3_mulDivCtrl_isSigned;
  reg                 entriesNext_3_mulDivCtrl_isWordOp;
  reg                 entryValidsNext_0;
  reg                 entryValidsNext_1;
  reg                 entryValidsNext_2;
  reg                 entryValidsNext_3;
  wire                when_IssueQueueComponent_l186;
  wire                when_IssueQueueComponent_l187;
  wire                when_IssueQueueComponent_l186_1;
  wire                when_IssueQueueComponent_l187_1;
  wire                when_IssueQueueComponent_l186_2;
  wire                when_IssueQueueComponent_l187_2;
  wire                when_IssueQueueComponent_l186_3;
  wire                when_IssueQueueComponent_l187_3;
  wire       [3:0]    _zz_1;
  wire                io_allocateIn_fire;
  wire       [3:0]    _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_entriesNext_0_src1Ready;
  wire                _zz_entriesNext_0_src2Ready;
  wire       [3:0]    _zz_7;
  wire                when_IssueQueueComponent_l212;
  wire                when_IssueQueueComponent_l215;
  wire                when_IssueQueueComponent_l212_1;
  wire                when_IssueQueueComponent_l215_1;
  wire                when_IssueQueueComponent_l212_2;
  wire                when_IssueQueueComponent_l215_2;
  wire                when_IssueQueueComponent_l212_3;
  wire                when_IssueQueueComponent_l215_3;
  wire                when_IssueQueueComponent_l212_4;
  wire                when_IssueQueueComponent_l215_4;
  wire       [2:0]    _zz_currentValidCount;
  wire       [2:0]    _zz_currentValidCount_1;
  wire       [2:0]    _zz_currentValidCount_2;
  wire       [2:0]    _zz_currentValidCount_3;
  wire       [2:0]    _zz_currentValidCount_4;
  wire       [2:0]    _zz_currentValidCount_5;
  wire       [2:0]    _zz_currentValidCount_6;
  wire       [2:0]    _zz_currentValidCount_7;
  wire       [2:0]    currentValidCount;
  wire                logCondition;
  wire                when_IssueQueueComponent_l256;
  `ifndef SYNTHESIS
  reg [87:0] io_allocateIn_payload_uop_decoded_uopCode_string;
  reg [151:0] io_allocateIn_payload_uop_decoded_exeUnit_string;
  reg [71:0] io_allocateIn_payload_uop_decoded_isa_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] io_allocateIn_payload_uop_decoded_immUsage_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] io_allocateIn_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_allocateIn_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] io_issueOut_payload_uop_decoded_uopCode_string;
  reg [151:0] io_issueOut_payload_uop_decoded_exeUnit_string;
  reg [71:0] io_issueOut_payload_uop_decoded_isa_string;
  reg [39:0] io_issueOut_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] io_issueOut_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] io_issueOut_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] io_issueOut_payload_uop_decoded_immUsage_string;
  reg [39:0] io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] io_issueOut_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] io_issueOut_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_issueOut_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] entries_0_uop_decoded_uopCode_string;
  reg [151:0] entries_0_uop_decoded_exeUnit_string;
  reg [71:0] entries_0_uop_decoded_isa_string;
  reg [39:0] entries_0_uop_decoded_archDest_rtype_string;
  reg [39:0] entries_0_uop_decoded_archSrc1_rtype_string;
  reg [39:0] entries_0_uop_decoded_archSrc2_rtype_string;
  reg [103:0] entries_0_uop_decoded_immUsage_string;
  reg [39:0] entries_0_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] entries_0_uop_decoded_memCtrl_size_string;
  reg [87:0] entries_0_uop_decoded_branchCtrl_condition_string;
  reg [39:0] entries_0_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] entries_0_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] entries_0_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] entries_0_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] entries_0_uop_decoded_decodeExceptionCode_string;
  reg [87:0] entries_1_uop_decoded_uopCode_string;
  reg [151:0] entries_1_uop_decoded_exeUnit_string;
  reg [71:0] entries_1_uop_decoded_isa_string;
  reg [39:0] entries_1_uop_decoded_archDest_rtype_string;
  reg [39:0] entries_1_uop_decoded_archSrc1_rtype_string;
  reg [39:0] entries_1_uop_decoded_archSrc2_rtype_string;
  reg [103:0] entries_1_uop_decoded_immUsage_string;
  reg [39:0] entries_1_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] entries_1_uop_decoded_memCtrl_size_string;
  reg [87:0] entries_1_uop_decoded_branchCtrl_condition_string;
  reg [39:0] entries_1_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] entries_1_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] entries_1_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] entries_1_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] entries_1_uop_decoded_decodeExceptionCode_string;
  reg [87:0] entries_2_uop_decoded_uopCode_string;
  reg [151:0] entries_2_uop_decoded_exeUnit_string;
  reg [71:0] entries_2_uop_decoded_isa_string;
  reg [39:0] entries_2_uop_decoded_archDest_rtype_string;
  reg [39:0] entries_2_uop_decoded_archSrc1_rtype_string;
  reg [39:0] entries_2_uop_decoded_archSrc2_rtype_string;
  reg [103:0] entries_2_uop_decoded_immUsage_string;
  reg [39:0] entries_2_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] entries_2_uop_decoded_memCtrl_size_string;
  reg [87:0] entries_2_uop_decoded_branchCtrl_condition_string;
  reg [39:0] entries_2_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] entries_2_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] entries_2_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] entries_2_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] entries_2_uop_decoded_decodeExceptionCode_string;
  reg [87:0] entries_3_uop_decoded_uopCode_string;
  reg [151:0] entries_3_uop_decoded_exeUnit_string;
  reg [71:0] entries_3_uop_decoded_isa_string;
  reg [39:0] entries_3_uop_decoded_archDest_rtype_string;
  reg [39:0] entries_3_uop_decoded_archSrc1_rtype_string;
  reg [39:0] entries_3_uop_decoded_archSrc2_rtype_string;
  reg [103:0] entries_3_uop_decoded_immUsage_string;
  reg [39:0] entries_3_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] entries_3_uop_decoded_memCtrl_size_string;
  reg [87:0] entries_3_uop_decoded_branchCtrl_condition_string;
  reg [39:0] entries_3_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] entries_3_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] entries_3_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] entries_3_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] entries_3_uop_decoded_decodeExceptionCode_string;
  reg [87:0] _zz_io_issueOut_payload_uop_decoded_uopCode_string;
  reg [151:0] _zz_io_issueOut_payload_uop_decoded_exeUnit_string;
  reg [71:0] _zz_io_issueOut_payload_uop_decoded_isa_string;
  reg [39:0] _zz_io_issueOut_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] _zz_io_issueOut_payload_uop_decoded_immUsage_string;
  reg [39:0] _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] _zz_io_issueOut_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] entriesNext_0_uop_decoded_uopCode_string;
  reg [151:0] entriesNext_0_uop_decoded_exeUnit_string;
  reg [71:0] entriesNext_0_uop_decoded_isa_string;
  reg [39:0] entriesNext_0_uop_decoded_archDest_rtype_string;
  reg [39:0] entriesNext_0_uop_decoded_archSrc1_rtype_string;
  reg [39:0] entriesNext_0_uop_decoded_archSrc2_rtype_string;
  reg [103:0] entriesNext_0_uop_decoded_immUsage_string;
  reg [39:0] entriesNext_0_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] entriesNext_0_uop_decoded_memCtrl_size_string;
  reg [87:0] entriesNext_0_uop_decoded_branchCtrl_condition_string;
  reg [39:0] entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] entriesNext_0_uop_decoded_decodeExceptionCode_string;
  reg [87:0] entriesNext_1_uop_decoded_uopCode_string;
  reg [151:0] entriesNext_1_uop_decoded_exeUnit_string;
  reg [71:0] entriesNext_1_uop_decoded_isa_string;
  reg [39:0] entriesNext_1_uop_decoded_archDest_rtype_string;
  reg [39:0] entriesNext_1_uop_decoded_archSrc1_rtype_string;
  reg [39:0] entriesNext_1_uop_decoded_archSrc2_rtype_string;
  reg [103:0] entriesNext_1_uop_decoded_immUsage_string;
  reg [39:0] entriesNext_1_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] entriesNext_1_uop_decoded_memCtrl_size_string;
  reg [87:0] entriesNext_1_uop_decoded_branchCtrl_condition_string;
  reg [39:0] entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] entriesNext_1_uop_decoded_decodeExceptionCode_string;
  reg [87:0] entriesNext_2_uop_decoded_uopCode_string;
  reg [151:0] entriesNext_2_uop_decoded_exeUnit_string;
  reg [71:0] entriesNext_2_uop_decoded_isa_string;
  reg [39:0] entriesNext_2_uop_decoded_archDest_rtype_string;
  reg [39:0] entriesNext_2_uop_decoded_archSrc1_rtype_string;
  reg [39:0] entriesNext_2_uop_decoded_archSrc2_rtype_string;
  reg [103:0] entriesNext_2_uop_decoded_immUsage_string;
  reg [39:0] entriesNext_2_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] entriesNext_2_uop_decoded_memCtrl_size_string;
  reg [87:0] entriesNext_2_uop_decoded_branchCtrl_condition_string;
  reg [39:0] entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] entriesNext_2_uop_decoded_decodeExceptionCode_string;
  reg [87:0] entriesNext_3_uop_decoded_uopCode_string;
  reg [151:0] entriesNext_3_uop_decoded_exeUnit_string;
  reg [71:0] entriesNext_3_uop_decoded_isa_string;
  reg [39:0] entriesNext_3_uop_decoded_archDest_rtype_string;
  reg [39:0] entriesNext_3_uop_decoded_archSrc1_rtype_string;
  reg [39:0] entriesNext_3_uop_decoded_archSrc2_rtype_string;
  reg [103:0] entriesNext_3_uop_decoded_immUsage_string;
  reg [39:0] entriesNext_3_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] entriesNext_3_uop_decoded_memCtrl_size_string;
  reg [87:0] entriesNext_3_uop_decoded_branchCtrl_condition_string;
  reg [39:0] entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] entriesNext_3_uop_decoded_decodeExceptionCode_string;
  `endif


  assign _zz_issueRequestMask_ohFirst_masked = (issueRequestMask_ohFirst_input - 4'b0001);
  assign _zz_allocationMask_1 = (_zz_allocationMask - 4'b0001);
  assign _zz_currentValidCount_12 = entryValids_3;
  assign _zz_currentValidCount_11 = {2'd0, _zz_currentValidCount_12};
  assign _zz_currentValidCount_9 = {entryValids_2,{entryValids_1,entryValids_0}};
  always @(*) begin
    case(issueIdx)
      2'b00 : begin
        _zz__zz_io_issueOut_payload_uop_decoded_uopCode = entries_0_uop_decoded_uopCode;
        _zz__zz_io_issueOut_payload_uop_decoded_exeUnit = entries_0_uop_decoded_exeUnit;
        _zz__zz_io_issueOut_payload_uop_decoded_isa = entries_0_uop_decoded_isa;
        _zz__zz_io_issueOut_payload_uop_decoded_archDest_rtype = entries_0_uop_decoded_archDest_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_archSrc1_rtype = entries_0_uop_decoded_archSrc1_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_archSrc2_rtype = entries_0_uop_decoded_archSrc2_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_immUsage = entries_0_uop_decoded_immUsage;
        _zz__zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp = entries_0_uop_decoded_aluCtrl_logicOp;
        _zz__zz_io_issueOut_payload_uop_decoded_memCtrl_size = entries_0_uop_decoded_memCtrl_size;
        _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_condition = entries_0_uop_decoded_branchCtrl_condition;
        _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype = entries_0_uop_decoded_branchCtrl_linkReg_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = entries_0_uop_decoded_fpuCtrl_fpSizeSrc1;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = entries_0_uop_decoded_fpuCtrl_fpSizeSrc2;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest = entries_0_uop_decoded_fpuCtrl_fpSizeDest;
        _zz__zz_io_issueOut_payload_uop_decoded_decodeExceptionCode = entries_0_uop_decoded_decodeExceptionCode;
        _zz_io_issueOut_payload_uop_decoded_pc = entries_0_uop_decoded_pc;
        _zz_io_issueOut_payload_uop_decoded_isValid = entries_0_uop_decoded_isValid;
        _zz_io_issueOut_payload_uop_decoded_archDest_idx = entries_0_uop_decoded_archDest_idx;
        _zz_io_issueOut_payload_uop_decoded_writeArchDestEn = entries_0_uop_decoded_writeArchDestEn;
        _zz_io_issueOut_payload_uop_decoded_archSrc1_idx = entries_0_uop_decoded_archSrc1_idx;
        _zz_io_issueOut_payload_uop_decoded_useArchSrc1 = entries_0_uop_decoded_useArchSrc1;
        _zz_io_issueOut_payload_uop_decoded_archSrc2_idx = entries_0_uop_decoded_archSrc2_idx;
        _zz_io_issueOut_payload_uop_decoded_useArchSrc2 = entries_0_uop_decoded_useArchSrc2;
        _zz_io_issueOut_payload_uop_decoded_usePcForAddr = entries_0_uop_decoded_usePcForAddr;
        _zz_io_issueOut_payload_uop_decoded_imm = entries_0_uop_decoded_imm;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_valid = entries_0_uop_decoded_aluCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSub = entries_0_uop_decoded_aluCtrl_isSub;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isAdd = entries_0_uop_decoded_aluCtrl_isAdd;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSigned = entries_0_uop_decoded_aluCtrl_isSigned;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_valid = entries_0_uop_decoded_shiftCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRight = entries_0_uop_decoded_shiftCtrl_isRight;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic = entries_0_uop_decoded_shiftCtrl_isArithmetic;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate = entries_0_uop_decoded_shiftCtrl_isRotate;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord = entries_0_uop_decoded_shiftCtrl_isDoubleWord;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_valid = entries_0_uop_decoded_mulDivCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv = entries_0_uop_decoded_mulDivCtrl_isDiv;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned = entries_0_uop_decoded_mulDivCtrl_isSigned;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp = entries_0_uop_decoded_mulDivCtrl_isWordOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad = entries_0_uop_decoded_memCtrl_isSignedLoad;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isStore = entries_0_uop_decoded_memCtrl_isStore;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked = entries_0_uop_decoded_memCtrl_isLoadLinked;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond = entries_0_uop_decoded_memCtrl_isStoreCond;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_atomicOp = entries_0_uop_decoded_memCtrl_atomicOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isFence = entries_0_uop_decoded_memCtrl_isFence;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_fenceMode = entries_0_uop_decoded_memCtrl_fenceMode;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp = entries_0_uop_decoded_memCtrl_isCacheOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType = entries_0_uop_decoded_memCtrl_cacheOpType;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch = entries_0_uop_decoded_memCtrl_isPrefetch;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isJump = entries_0_uop_decoded_branchCtrl_isJump;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isLink = entries_0_uop_decoded_branchCtrl_isLink;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx = entries_0_uop_decoded_branchCtrl_linkReg_idx;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect = entries_0_uop_decoded_branchCtrl_isIndirect;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx = entries_0_uop_decoded_branchCtrl_laCfIdx;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_opType = entries_0_uop_decoded_fpuCtrl_opType;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode = entries_0_uop_decoded_fpuCtrl_roundingMode;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest = entries_0_uop_decoded_fpuCtrl_isIntegerDest;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt = entries_0_uop_decoded_fpuCtrl_isSignedCvt;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = entries_0_uop_decoded_fpuCtrl_fmaNegSrc1;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond = entries_0_uop_decoded_fpuCtrl_fcmpCond;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr = entries_0_uop_decoded_csrCtrl_csrAddr;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isWrite = entries_0_uop_decoded_csrCtrl_isWrite;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isRead = entries_0_uop_decoded_csrCtrl_isRead;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isExchange = entries_0_uop_decoded_csrCtrl_isExchange;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc = entries_0_uop_decoded_csrCtrl_useUimmAsSrc;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_sysCode = entries_0_uop_decoded_sysCtrl_sysCode;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn = entries_0_uop_decoded_sysCtrl_isExceptionReturn;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp = entries_0_uop_decoded_sysCtrl_isTlbOp;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType = entries_0_uop_decoded_sysCtrl_tlbOpType;
        _zz_io_issueOut_payload_uop_decoded_hasDecodeException = entries_0_uop_decoded_hasDecodeException;
        _zz_io_issueOut_payload_uop_decoded_isMicrocode = entries_0_uop_decoded_isMicrocode;
        _zz_io_issueOut_payload_uop_decoded_microcodeEntry = entries_0_uop_decoded_microcodeEntry;
        _zz_io_issueOut_payload_uop_decoded_isSerializing = entries_0_uop_decoded_isSerializing;
        _zz_io_issueOut_payload_uop_decoded_isBranchOrJump = entries_0_uop_decoded_isBranchOrJump;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_isTaken = entries_0_uop_decoded_branchPrediction_isTaken;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_target = entries_0_uop_decoded_branchPrediction_target;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted = entries_0_uop_decoded_branchPrediction_wasPredicted;
        _zz_io_issueOut_payload_uop_rename_physSrc1_idx = entries_0_uop_rename_physSrc1_idx;
        _zz_io_issueOut_payload_uop_rename_physSrc1IsFpr = entries_0_uop_rename_physSrc1IsFpr;
        _zz_io_issueOut_payload_uop_rename_physSrc2_idx = entries_0_uop_rename_physSrc2_idx;
        _zz_io_issueOut_payload_uop_rename_physSrc2IsFpr = entries_0_uop_rename_physSrc2IsFpr;
        _zz_io_issueOut_payload_uop_rename_physDest_idx = entries_0_uop_rename_physDest_idx;
        _zz_io_issueOut_payload_uop_rename_physDestIsFpr = entries_0_uop_rename_physDestIsFpr;
        _zz_io_issueOut_payload_uop_rename_oldPhysDest_idx = entries_0_uop_rename_oldPhysDest_idx;
        _zz_io_issueOut_payload_uop_rename_oldPhysDestIsFpr = entries_0_uop_rename_oldPhysDestIsFpr;
        _zz_io_issueOut_payload_uop_rename_allocatesPhysDest = entries_0_uop_rename_allocatesPhysDest;
        _zz_io_issueOut_payload_uop_rename_writesToPhysReg = entries_0_uop_rename_writesToPhysReg;
        _zz_io_issueOut_payload_uop_robPtr = entries_0_uop_robPtr;
        _zz_io_issueOut_payload_uop_uniqueId = entries_0_uop_uniqueId;
        _zz_io_issueOut_payload_uop_dispatched = entries_0_uop_dispatched;
        _zz_io_issueOut_payload_uop_executed = entries_0_uop_executed;
        _zz_io_issueOut_payload_uop_hasException = entries_0_uop_hasException;
        _zz_io_issueOut_payload_uop_exceptionCode = entries_0_uop_exceptionCode;
        _zz_io_issueOut_payload_robPtr = entries_0_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_0_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_0_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_0_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_0_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_0_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_0_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_0_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_0_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_0_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_0_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_0_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_0_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_0_src2IsFpr;
        _zz_io_issueOut_payload_mulDivCtrl_valid = entries_0_mulDivCtrl_valid;
        _zz_io_issueOut_payload_mulDivCtrl_isDiv = entries_0_mulDivCtrl_isDiv;
        _zz_io_issueOut_payload_mulDivCtrl_isSigned = entries_0_mulDivCtrl_isSigned;
        _zz_io_issueOut_payload_mulDivCtrl_isWordOp = entries_0_mulDivCtrl_isWordOp;
      end
      2'b01 : begin
        _zz__zz_io_issueOut_payload_uop_decoded_uopCode = entries_1_uop_decoded_uopCode;
        _zz__zz_io_issueOut_payload_uop_decoded_exeUnit = entries_1_uop_decoded_exeUnit;
        _zz__zz_io_issueOut_payload_uop_decoded_isa = entries_1_uop_decoded_isa;
        _zz__zz_io_issueOut_payload_uop_decoded_archDest_rtype = entries_1_uop_decoded_archDest_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_archSrc1_rtype = entries_1_uop_decoded_archSrc1_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_archSrc2_rtype = entries_1_uop_decoded_archSrc2_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_immUsage = entries_1_uop_decoded_immUsage;
        _zz__zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp = entries_1_uop_decoded_aluCtrl_logicOp;
        _zz__zz_io_issueOut_payload_uop_decoded_memCtrl_size = entries_1_uop_decoded_memCtrl_size;
        _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_condition = entries_1_uop_decoded_branchCtrl_condition;
        _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype = entries_1_uop_decoded_branchCtrl_linkReg_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = entries_1_uop_decoded_fpuCtrl_fpSizeSrc1;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = entries_1_uop_decoded_fpuCtrl_fpSizeSrc2;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest = entries_1_uop_decoded_fpuCtrl_fpSizeDest;
        _zz__zz_io_issueOut_payload_uop_decoded_decodeExceptionCode = entries_1_uop_decoded_decodeExceptionCode;
        _zz_io_issueOut_payload_uop_decoded_pc = entries_1_uop_decoded_pc;
        _zz_io_issueOut_payload_uop_decoded_isValid = entries_1_uop_decoded_isValid;
        _zz_io_issueOut_payload_uop_decoded_archDest_idx = entries_1_uop_decoded_archDest_idx;
        _zz_io_issueOut_payload_uop_decoded_writeArchDestEn = entries_1_uop_decoded_writeArchDestEn;
        _zz_io_issueOut_payload_uop_decoded_archSrc1_idx = entries_1_uop_decoded_archSrc1_idx;
        _zz_io_issueOut_payload_uop_decoded_useArchSrc1 = entries_1_uop_decoded_useArchSrc1;
        _zz_io_issueOut_payload_uop_decoded_archSrc2_idx = entries_1_uop_decoded_archSrc2_idx;
        _zz_io_issueOut_payload_uop_decoded_useArchSrc2 = entries_1_uop_decoded_useArchSrc2;
        _zz_io_issueOut_payload_uop_decoded_usePcForAddr = entries_1_uop_decoded_usePcForAddr;
        _zz_io_issueOut_payload_uop_decoded_imm = entries_1_uop_decoded_imm;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_valid = entries_1_uop_decoded_aluCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSub = entries_1_uop_decoded_aluCtrl_isSub;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isAdd = entries_1_uop_decoded_aluCtrl_isAdd;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSigned = entries_1_uop_decoded_aluCtrl_isSigned;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_valid = entries_1_uop_decoded_shiftCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRight = entries_1_uop_decoded_shiftCtrl_isRight;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic = entries_1_uop_decoded_shiftCtrl_isArithmetic;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate = entries_1_uop_decoded_shiftCtrl_isRotate;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord = entries_1_uop_decoded_shiftCtrl_isDoubleWord;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_valid = entries_1_uop_decoded_mulDivCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv = entries_1_uop_decoded_mulDivCtrl_isDiv;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned = entries_1_uop_decoded_mulDivCtrl_isSigned;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp = entries_1_uop_decoded_mulDivCtrl_isWordOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad = entries_1_uop_decoded_memCtrl_isSignedLoad;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isStore = entries_1_uop_decoded_memCtrl_isStore;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked = entries_1_uop_decoded_memCtrl_isLoadLinked;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond = entries_1_uop_decoded_memCtrl_isStoreCond;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_atomicOp = entries_1_uop_decoded_memCtrl_atomicOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isFence = entries_1_uop_decoded_memCtrl_isFence;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_fenceMode = entries_1_uop_decoded_memCtrl_fenceMode;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp = entries_1_uop_decoded_memCtrl_isCacheOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType = entries_1_uop_decoded_memCtrl_cacheOpType;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch = entries_1_uop_decoded_memCtrl_isPrefetch;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isJump = entries_1_uop_decoded_branchCtrl_isJump;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isLink = entries_1_uop_decoded_branchCtrl_isLink;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx = entries_1_uop_decoded_branchCtrl_linkReg_idx;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect = entries_1_uop_decoded_branchCtrl_isIndirect;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx = entries_1_uop_decoded_branchCtrl_laCfIdx;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_opType = entries_1_uop_decoded_fpuCtrl_opType;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode = entries_1_uop_decoded_fpuCtrl_roundingMode;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest = entries_1_uop_decoded_fpuCtrl_isIntegerDest;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt = entries_1_uop_decoded_fpuCtrl_isSignedCvt;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = entries_1_uop_decoded_fpuCtrl_fmaNegSrc1;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond = entries_1_uop_decoded_fpuCtrl_fcmpCond;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr = entries_1_uop_decoded_csrCtrl_csrAddr;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isWrite = entries_1_uop_decoded_csrCtrl_isWrite;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isRead = entries_1_uop_decoded_csrCtrl_isRead;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isExchange = entries_1_uop_decoded_csrCtrl_isExchange;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc = entries_1_uop_decoded_csrCtrl_useUimmAsSrc;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_sysCode = entries_1_uop_decoded_sysCtrl_sysCode;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn = entries_1_uop_decoded_sysCtrl_isExceptionReturn;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp = entries_1_uop_decoded_sysCtrl_isTlbOp;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType = entries_1_uop_decoded_sysCtrl_tlbOpType;
        _zz_io_issueOut_payload_uop_decoded_hasDecodeException = entries_1_uop_decoded_hasDecodeException;
        _zz_io_issueOut_payload_uop_decoded_isMicrocode = entries_1_uop_decoded_isMicrocode;
        _zz_io_issueOut_payload_uop_decoded_microcodeEntry = entries_1_uop_decoded_microcodeEntry;
        _zz_io_issueOut_payload_uop_decoded_isSerializing = entries_1_uop_decoded_isSerializing;
        _zz_io_issueOut_payload_uop_decoded_isBranchOrJump = entries_1_uop_decoded_isBranchOrJump;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_isTaken = entries_1_uop_decoded_branchPrediction_isTaken;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_target = entries_1_uop_decoded_branchPrediction_target;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted = entries_1_uop_decoded_branchPrediction_wasPredicted;
        _zz_io_issueOut_payload_uop_rename_physSrc1_idx = entries_1_uop_rename_physSrc1_idx;
        _zz_io_issueOut_payload_uop_rename_physSrc1IsFpr = entries_1_uop_rename_physSrc1IsFpr;
        _zz_io_issueOut_payload_uop_rename_physSrc2_idx = entries_1_uop_rename_physSrc2_idx;
        _zz_io_issueOut_payload_uop_rename_physSrc2IsFpr = entries_1_uop_rename_physSrc2IsFpr;
        _zz_io_issueOut_payload_uop_rename_physDest_idx = entries_1_uop_rename_physDest_idx;
        _zz_io_issueOut_payload_uop_rename_physDestIsFpr = entries_1_uop_rename_physDestIsFpr;
        _zz_io_issueOut_payload_uop_rename_oldPhysDest_idx = entries_1_uop_rename_oldPhysDest_idx;
        _zz_io_issueOut_payload_uop_rename_oldPhysDestIsFpr = entries_1_uop_rename_oldPhysDestIsFpr;
        _zz_io_issueOut_payload_uop_rename_allocatesPhysDest = entries_1_uop_rename_allocatesPhysDest;
        _zz_io_issueOut_payload_uop_rename_writesToPhysReg = entries_1_uop_rename_writesToPhysReg;
        _zz_io_issueOut_payload_uop_robPtr = entries_1_uop_robPtr;
        _zz_io_issueOut_payload_uop_uniqueId = entries_1_uop_uniqueId;
        _zz_io_issueOut_payload_uop_dispatched = entries_1_uop_dispatched;
        _zz_io_issueOut_payload_uop_executed = entries_1_uop_executed;
        _zz_io_issueOut_payload_uop_hasException = entries_1_uop_hasException;
        _zz_io_issueOut_payload_uop_exceptionCode = entries_1_uop_exceptionCode;
        _zz_io_issueOut_payload_robPtr = entries_1_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_1_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_1_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_1_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_1_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_1_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_1_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_1_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_1_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_1_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_1_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_1_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_1_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_1_src2IsFpr;
        _zz_io_issueOut_payload_mulDivCtrl_valid = entries_1_mulDivCtrl_valid;
        _zz_io_issueOut_payload_mulDivCtrl_isDiv = entries_1_mulDivCtrl_isDiv;
        _zz_io_issueOut_payload_mulDivCtrl_isSigned = entries_1_mulDivCtrl_isSigned;
        _zz_io_issueOut_payload_mulDivCtrl_isWordOp = entries_1_mulDivCtrl_isWordOp;
      end
      2'b10 : begin
        _zz__zz_io_issueOut_payload_uop_decoded_uopCode = entries_2_uop_decoded_uopCode;
        _zz__zz_io_issueOut_payload_uop_decoded_exeUnit = entries_2_uop_decoded_exeUnit;
        _zz__zz_io_issueOut_payload_uop_decoded_isa = entries_2_uop_decoded_isa;
        _zz__zz_io_issueOut_payload_uop_decoded_archDest_rtype = entries_2_uop_decoded_archDest_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_archSrc1_rtype = entries_2_uop_decoded_archSrc1_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_archSrc2_rtype = entries_2_uop_decoded_archSrc2_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_immUsage = entries_2_uop_decoded_immUsage;
        _zz__zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp = entries_2_uop_decoded_aluCtrl_logicOp;
        _zz__zz_io_issueOut_payload_uop_decoded_memCtrl_size = entries_2_uop_decoded_memCtrl_size;
        _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_condition = entries_2_uop_decoded_branchCtrl_condition;
        _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype = entries_2_uop_decoded_branchCtrl_linkReg_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = entries_2_uop_decoded_fpuCtrl_fpSizeSrc1;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = entries_2_uop_decoded_fpuCtrl_fpSizeSrc2;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest = entries_2_uop_decoded_fpuCtrl_fpSizeDest;
        _zz__zz_io_issueOut_payload_uop_decoded_decodeExceptionCode = entries_2_uop_decoded_decodeExceptionCode;
        _zz_io_issueOut_payload_uop_decoded_pc = entries_2_uop_decoded_pc;
        _zz_io_issueOut_payload_uop_decoded_isValid = entries_2_uop_decoded_isValid;
        _zz_io_issueOut_payload_uop_decoded_archDest_idx = entries_2_uop_decoded_archDest_idx;
        _zz_io_issueOut_payload_uop_decoded_writeArchDestEn = entries_2_uop_decoded_writeArchDestEn;
        _zz_io_issueOut_payload_uop_decoded_archSrc1_idx = entries_2_uop_decoded_archSrc1_idx;
        _zz_io_issueOut_payload_uop_decoded_useArchSrc1 = entries_2_uop_decoded_useArchSrc1;
        _zz_io_issueOut_payload_uop_decoded_archSrc2_idx = entries_2_uop_decoded_archSrc2_idx;
        _zz_io_issueOut_payload_uop_decoded_useArchSrc2 = entries_2_uop_decoded_useArchSrc2;
        _zz_io_issueOut_payload_uop_decoded_usePcForAddr = entries_2_uop_decoded_usePcForAddr;
        _zz_io_issueOut_payload_uop_decoded_imm = entries_2_uop_decoded_imm;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_valid = entries_2_uop_decoded_aluCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSub = entries_2_uop_decoded_aluCtrl_isSub;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isAdd = entries_2_uop_decoded_aluCtrl_isAdd;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSigned = entries_2_uop_decoded_aluCtrl_isSigned;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_valid = entries_2_uop_decoded_shiftCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRight = entries_2_uop_decoded_shiftCtrl_isRight;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic = entries_2_uop_decoded_shiftCtrl_isArithmetic;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate = entries_2_uop_decoded_shiftCtrl_isRotate;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord = entries_2_uop_decoded_shiftCtrl_isDoubleWord;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_valid = entries_2_uop_decoded_mulDivCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv = entries_2_uop_decoded_mulDivCtrl_isDiv;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned = entries_2_uop_decoded_mulDivCtrl_isSigned;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp = entries_2_uop_decoded_mulDivCtrl_isWordOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad = entries_2_uop_decoded_memCtrl_isSignedLoad;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isStore = entries_2_uop_decoded_memCtrl_isStore;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked = entries_2_uop_decoded_memCtrl_isLoadLinked;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond = entries_2_uop_decoded_memCtrl_isStoreCond;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_atomicOp = entries_2_uop_decoded_memCtrl_atomicOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isFence = entries_2_uop_decoded_memCtrl_isFence;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_fenceMode = entries_2_uop_decoded_memCtrl_fenceMode;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp = entries_2_uop_decoded_memCtrl_isCacheOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType = entries_2_uop_decoded_memCtrl_cacheOpType;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch = entries_2_uop_decoded_memCtrl_isPrefetch;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isJump = entries_2_uop_decoded_branchCtrl_isJump;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isLink = entries_2_uop_decoded_branchCtrl_isLink;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx = entries_2_uop_decoded_branchCtrl_linkReg_idx;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect = entries_2_uop_decoded_branchCtrl_isIndirect;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx = entries_2_uop_decoded_branchCtrl_laCfIdx;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_opType = entries_2_uop_decoded_fpuCtrl_opType;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode = entries_2_uop_decoded_fpuCtrl_roundingMode;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest = entries_2_uop_decoded_fpuCtrl_isIntegerDest;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt = entries_2_uop_decoded_fpuCtrl_isSignedCvt;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = entries_2_uop_decoded_fpuCtrl_fmaNegSrc1;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond = entries_2_uop_decoded_fpuCtrl_fcmpCond;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr = entries_2_uop_decoded_csrCtrl_csrAddr;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isWrite = entries_2_uop_decoded_csrCtrl_isWrite;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isRead = entries_2_uop_decoded_csrCtrl_isRead;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isExchange = entries_2_uop_decoded_csrCtrl_isExchange;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc = entries_2_uop_decoded_csrCtrl_useUimmAsSrc;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_sysCode = entries_2_uop_decoded_sysCtrl_sysCode;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn = entries_2_uop_decoded_sysCtrl_isExceptionReturn;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp = entries_2_uop_decoded_sysCtrl_isTlbOp;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType = entries_2_uop_decoded_sysCtrl_tlbOpType;
        _zz_io_issueOut_payload_uop_decoded_hasDecodeException = entries_2_uop_decoded_hasDecodeException;
        _zz_io_issueOut_payload_uop_decoded_isMicrocode = entries_2_uop_decoded_isMicrocode;
        _zz_io_issueOut_payload_uop_decoded_microcodeEntry = entries_2_uop_decoded_microcodeEntry;
        _zz_io_issueOut_payload_uop_decoded_isSerializing = entries_2_uop_decoded_isSerializing;
        _zz_io_issueOut_payload_uop_decoded_isBranchOrJump = entries_2_uop_decoded_isBranchOrJump;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_isTaken = entries_2_uop_decoded_branchPrediction_isTaken;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_target = entries_2_uop_decoded_branchPrediction_target;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted = entries_2_uop_decoded_branchPrediction_wasPredicted;
        _zz_io_issueOut_payload_uop_rename_physSrc1_idx = entries_2_uop_rename_physSrc1_idx;
        _zz_io_issueOut_payload_uop_rename_physSrc1IsFpr = entries_2_uop_rename_physSrc1IsFpr;
        _zz_io_issueOut_payload_uop_rename_physSrc2_idx = entries_2_uop_rename_physSrc2_idx;
        _zz_io_issueOut_payload_uop_rename_physSrc2IsFpr = entries_2_uop_rename_physSrc2IsFpr;
        _zz_io_issueOut_payload_uop_rename_physDest_idx = entries_2_uop_rename_physDest_idx;
        _zz_io_issueOut_payload_uop_rename_physDestIsFpr = entries_2_uop_rename_physDestIsFpr;
        _zz_io_issueOut_payload_uop_rename_oldPhysDest_idx = entries_2_uop_rename_oldPhysDest_idx;
        _zz_io_issueOut_payload_uop_rename_oldPhysDestIsFpr = entries_2_uop_rename_oldPhysDestIsFpr;
        _zz_io_issueOut_payload_uop_rename_allocatesPhysDest = entries_2_uop_rename_allocatesPhysDest;
        _zz_io_issueOut_payload_uop_rename_writesToPhysReg = entries_2_uop_rename_writesToPhysReg;
        _zz_io_issueOut_payload_uop_robPtr = entries_2_uop_robPtr;
        _zz_io_issueOut_payload_uop_uniqueId = entries_2_uop_uniqueId;
        _zz_io_issueOut_payload_uop_dispatched = entries_2_uop_dispatched;
        _zz_io_issueOut_payload_uop_executed = entries_2_uop_executed;
        _zz_io_issueOut_payload_uop_hasException = entries_2_uop_hasException;
        _zz_io_issueOut_payload_uop_exceptionCode = entries_2_uop_exceptionCode;
        _zz_io_issueOut_payload_robPtr = entries_2_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_2_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_2_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_2_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_2_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_2_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_2_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_2_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_2_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_2_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_2_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_2_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_2_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_2_src2IsFpr;
        _zz_io_issueOut_payload_mulDivCtrl_valid = entries_2_mulDivCtrl_valid;
        _zz_io_issueOut_payload_mulDivCtrl_isDiv = entries_2_mulDivCtrl_isDiv;
        _zz_io_issueOut_payload_mulDivCtrl_isSigned = entries_2_mulDivCtrl_isSigned;
        _zz_io_issueOut_payload_mulDivCtrl_isWordOp = entries_2_mulDivCtrl_isWordOp;
      end
      default : begin
        _zz__zz_io_issueOut_payload_uop_decoded_uopCode = entries_3_uop_decoded_uopCode;
        _zz__zz_io_issueOut_payload_uop_decoded_exeUnit = entries_3_uop_decoded_exeUnit;
        _zz__zz_io_issueOut_payload_uop_decoded_isa = entries_3_uop_decoded_isa;
        _zz__zz_io_issueOut_payload_uop_decoded_archDest_rtype = entries_3_uop_decoded_archDest_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_archSrc1_rtype = entries_3_uop_decoded_archSrc1_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_archSrc2_rtype = entries_3_uop_decoded_archSrc2_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_immUsage = entries_3_uop_decoded_immUsage;
        _zz__zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp = entries_3_uop_decoded_aluCtrl_logicOp;
        _zz__zz_io_issueOut_payload_uop_decoded_memCtrl_size = entries_3_uop_decoded_memCtrl_size;
        _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_condition = entries_3_uop_decoded_branchCtrl_condition;
        _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype = entries_3_uop_decoded_branchCtrl_linkReg_rtype;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = entries_3_uop_decoded_fpuCtrl_fpSizeSrc1;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = entries_3_uop_decoded_fpuCtrl_fpSizeSrc2;
        _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest = entries_3_uop_decoded_fpuCtrl_fpSizeDest;
        _zz__zz_io_issueOut_payload_uop_decoded_decodeExceptionCode = entries_3_uop_decoded_decodeExceptionCode;
        _zz_io_issueOut_payload_uop_decoded_pc = entries_3_uop_decoded_pc;
        _zz_io_issueOut_payload_uop_decoded_isValid = entries_3_uop_decoded_isValid;
        _zz_io_issueOut_payload_uop_decoded_archDest_idx = entries_3_uop_decoded_archDest_idx;
        _zz_io_issueOut_payload_uop_decoded_writeArchDestEn = entries_3_uop_decoded_writeArchDestEn;
        _zz_io_issueOut_payload_uop_decoded_archSrc1_idx = entries_3_uop_decoded_archSrc1_idx;
        _zz_io_issueOut_payload_uop_decoded_useArchSrc1 = entries_3_uop_decoded_useArchSrc1;
        _zz_io_issueOut_payload_uop_decoded_archSrc2_idx = entries_3_uop_decoded_archSrc2_idx;
        _zz_io_issueOut_payload_uop_decoded_useArchSrc2 = entries_3_uop_decoded_useArchSrc2;
        _zz_io_issueOut_payload_uop_decoded_usePcForAddr = entries_3_uop_decoded_usePcForAddr;
        _zz_io_issueOut_payload_uop_decoded_imm = entries_3_uop_decoded_imm;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_valid = entries_3_uop_decoded_aluCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSub = entries_3_uop_decoded_aluCtrl_isSub;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isAdd = entries_3_uop_decoded_aluCtrl_isAdd;
        _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSigned = entries_3_uop_decoded_aluCtrl_isSigned;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_valid = entries_3_uop_decoded_shiftCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRight = entries_3_uop_decoded_shiftCtrl_isRight;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic = entries_3_uop_decoded_shiftCtrl_isArithmetic;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate = entries_3_uop_decoded_shiftCtrl_isRotate;
        _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord = entries_3_uop_decoded_shiftCtrl_isDoubleWord;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_valid = entries_3_uop_decoded_mulDivCtrl_valid;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv = entries_3_uop_decoded_mulDivCtrl_isDiv;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned = entries_3_uop_decoded_mulDivCtrl_isSigned;
        _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp = entries_3_uop_decoded_mulDivCtrl_isWordOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad = entries_3_uop_decoded_memCtrl_isSignedLoad;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isStore = entries_3_uop_decoded_memCtrl_isStore;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked = entries_3_uop_decoded_memCtrl_isLoadLinked;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond = entries_3_uop_decoded_memCtrl_isStoreCond;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_atomicOp = entries_3_uop_decoded_memCtrl_atomicOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isFence = entries_3_uop_decoded_memCtrl_isFence;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_fenceMode = entries_3_uop_decoded_memCtrl_fenceMode;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp = entries_3_uop_decoded_memCtrl_isCacheOp;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType = entries_3_uop_decoded_memCtrl_cacheOpType;
        _zz_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch = entries_3_uop_decoded_memCtrl_isPrefetch;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isJump = entries_3_uop_decoded_branchCtrl_isJump;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isLink = entries_3_uop_decoded_branchCtrl_isLink;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx = entries_3_uop_decoded_branchCtrl_linkReg_idx;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect = entries_3_uop_decoded_branchCtrl_isIndirect;
        _zz_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx = entries_3_uop_decoded_branchCtrl_laCfIdx;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_opType = entries_3_uop_decoded_fpuCtrl_opType;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode = entries_3_uop_decoded_fpuCtrl_roundingMode;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest = entries_3_uop_decoded_fpuCtrl_isIntegerDest;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt = entries_3_uop_decoded_fpuCtrl_isSignedCvt;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = entries_3_uop_decoded_fpuCtrl_fmaNegSrc1;
        _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond = entries_3_uop_decoded_fpuCtrl_fcmpCond;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr = entries_3_uop_decoded_csrCtrl_csrAddr;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isWrite = entries_3_uop_decoded_csrCtrl_isWrite;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isRead = entries_3_uop_decoded_csrCtrl_isRead;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_isExchange = entries_3_uop_decoded_csrCtrl_isExchange;
        _zz_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc = entries_3_uop_decoded_csrCtrl_useUimmAsSrc;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_sysCode = entries_3_uop_decoded_sysCtrl_sysCode;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn = entries_3_uop_decoded_sysCtrl_isExceptionReturn;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp = entries_3_uop_decoded_sysCtrl_isTlbOp;
        _zz_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType = entries_3_uop_decoded_sysCtrl_tlbOpType;
        _zz_io_issueOut_payload_uop_decoded_hasDecodeException = entries_3_uop_decoded_hasDecodeException;
        _zz_io_issueOut_payload_uop_decoded_isMicrocode = entries_3_uop_decoded_isMicrocode;
        _zz_io_issueOut_payload_uop_decoded_microcodeEntry = entries_3_uop_decoded_microcodeEntry;
        _zz_io_issueOut_payload_uop_decoded_isSerializing = entries_3_uop_decoded_isSerializing;
        _zz_io_issueOut_payload_uop_decoded_isBranchOrJump = entries_3_uop_decoded_isBranchOrJump;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_isTaken = entries_3_uop_decoded_branchPrediction_isTaken;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_target = entries_3_uop_decoded_branchPrediction_target;
        _zz_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted = entries_3_uop_decoded_branchPrediction_wasPredicted;
        _zz_io_issueOut_payload_uop_rename_physSrc1_idx = entries_3_uop_rename_physSrc1_idx;
        _zz_io_issueOut_payload_uop_rename_physSrc1IsFpr = entries_3_uop_rename_physSrc1IsFpr;
        _zz_io_issueOut_payload_uop_rename_physSrc2_idx = entries_3_uop_rename_physSrc2_idx;
        _zz_io_issueOut_payload_uop_rename_physSrc2IsFpr = entries_3_uop_rename_physSrc2IsFpr;
        _zz_io_issueOut_payload_uop_rename_physDest_idx = entries_3_uop_rename_physDest_idx;
        _zz_io_issueOut_payload_uop_rename_physDestIsFpr = entries_3_uop_rename_physDestIsFpr;
        _zz_io_issueOut_payload_uop_rename_oldPhysDest_idx = entries_3_uop_rename_oldPhysDest_idx;
        _zz_io_issueOut_payload_uop_rename_oldPhysDestIsFpr = entries_3_uop_rename_oldPhysDestIsFpr;
        _zz_io_issueOut_payload_uop_rename_allocatesPhysDest = entries_3_uop_rename_allocatesPhysDest;
        _zz_io_issueOut_payload_uop_rename_writesToPhysReg = entries_3_uop_rename_writesToPhysReg;
        _zz_io_issueOut_payload_uop_robPtr = entries_3_uop_robPtr;
        _zz_io_issueOut_payload_uop_uniqueId = entries_3_uop_uniqueId;
        _zz_io_issueOut_payload_uop_dispatched = entries_3_uop_dispatched;
        _zz_io_issueOut_payload_uop_executed = entries_3_uop_executed;
        _zz_io_issueOut_payload_uop_hasException = entries_3_uop_hasException;
        _zz_io_issueOut_payload_uop_exceptionCode = entries_3_uop_exceptionCode;
        _zz_io_issueOut_payload_robPtr = entries_3_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_3_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_3_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_3_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_3_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_3_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_3_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_3_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_3_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_3_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_3_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_3_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_3_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_3_src2IsFpr;
        _zz_io_issueOut_payload_mulDivCtrl_valid = entries_3_mulDivCtrl_valid;
        _zz_io_issueOut_payload_mulDivCtrl_isDiv = entries_3_mulDivCtrl_isDiv;
        _zz_io_issueOut_payload_mulDivCtrl_isSigned = entries_3_mulDivCtrl_isSigned;
        _zz_io_issueOut_payload_mulDivCtrl_isWordOp = entries_3_mulDivCtrl_isWordOp;
      end
    endcase
  end

  always @(*) begin
    case(_zz_currentValidCount_9)
      3'b000 : _zz_currentValidCount_8 = _zz_currentValidCount;
      3'b001 : _zz_currentValidCount_8 = _zz_currentValidCount_1;
      3'b010 : _zz_currentValidCount_8 = _zz_currentValidCount_2;
      3'b011 : _zz_currentValidCount_8 = _zz_currentValidCount_3;
      3'b100 : _zz_currentValidCount_8 = _zz_currentValidCount_4;
      3'b101 : _zz_currentValidCount_8 = _zz_currentValidCount_5;
      3'b110 : _zz_currentValidCount_8 = _zz_currentValidCount_6;
      default : _zz_currentValidCount_8 = _zz_currentValidCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_currentValidCount_11)
      3'b000 : _zz_currentValidCount_10 = _zz_currentValidCount;
      3'b001 : _zz_currentValidCount_10 = _zz_currentValidCount_1;
      3'b010 : _zz_currentValidCount_10 = _zz_currentValidCount_2;
      3'b011 : _zz_currentValidCount_10 = _zz_currentValidCount_3;
      3'b100 : _zz_currentValidCount_10 = _zz_currentValidCount_4;
      3'b101 : _zz_currentValidCount_10 = _zz_currentValidCount_5;
      3'b110 : _zz_currentValidCount_10 = _zz_currentValidCount_6;
      default : _zz_currentValidCount_10 = _zz_currentValidCount_7;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : io_allocateIn_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_allocateIn_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_allocateIn_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_allocateIn_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_allocateIn_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_allocateIn_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_allocateIn_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_allocateIn_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_allocateIn_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_allocateIn_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_allocateIn_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_allocateIn_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_allocateIn_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_allocateIn_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_allocateIn_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_allocateIn_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_allocateIn_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : io_allocateIn_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : io_allocateIn_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_allocateIn_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_allocateIn_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_allocateIn_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_allocateIn_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_allocateIn_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_allocateIn_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_isa)
      IsaType_UNKNOWN : io_allocateIn_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_allocateIn_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : io_allocateIn_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_allocateIn_payload_uop_decoded_isa_string = "LOONGARCH";
      default : io_allocateIn_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : io_allocateIn_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : io_allocateIn_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "D";
      default : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : io_issueOut_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_issueOut_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_issueOut_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_issueOut_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_issueOut_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_issueOut_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_issueOut_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_issueOut_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_issueOut_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_issueOut_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_issueOut_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_issueOut_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_issueOut_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_issueOut_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_issueOut_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_issueOut_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_issueOut_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_issueOut_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_issueOut_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_issueOut_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_issueOut_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_issueOut_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_issueOut_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_issueOut_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : io_issueOut_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : io_issueOut_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_issueOut_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_issueOut_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_issueOut_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_issueOut_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_issueOut_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_issueOut_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_issueOut_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_issueOut_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_issueOut_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_isa)
      IsaType_UNKNOWN : io_issueOut_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_issueOut_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : io_issueOut_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_issueOut_payload_uop_decoded_isa_string = "LOONGARCH";
      default : io_issueOut_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : io_issueOut_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_issueOut_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_issueOut_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_issueOut_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : io_issueOut_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : io_issueOut_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_issueOut_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_issueOut_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_issueOut_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_issueOut_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_issueOut_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_issueOut_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : io_issueOut_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : io_issueOut_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : io_issueOut_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : io_issueOut_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : io_issueOut_payload_uop_decoded_memCtrl_size_string = "D";
      default : io_issueOut_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_uopCode)
      BaseUopCode_NOP : entries_0_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : entries_0_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : entries_0_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : entries_0_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : entries_0_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : entries_0_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : entries_0_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : entries_0_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : entries_0_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : entries_0_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : entries_0_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : entries_0_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : entries_0_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : entries_0_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : entries_0_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : entries_0_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : entries_0_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : entries_0_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : entries_0_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : entries_0_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : entries_0_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : entries_0_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : entries_0_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : entries_0_uop_decoded_uopCode_string = "IDLE       ";
      default : entries_0_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_exeUnit)
      ExeUnitType_NONE : entries_0_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : entries_0_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : entries_0_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : entries_0_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : entries_0_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : entries_0_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : entries_0_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : entries_0_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : entries_0_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : entries_0_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_isa)
      IsaType_UNKNOWN : entries_0_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : entries_0_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : entries_0_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : entries_0_uop_decoded_isa_string = "LOONGARCH";
      default : entries_0_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_archDest_rtype)
      ArchRegType_GPR : entries_0_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_0_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_0_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_0_uop_decoded_archDest_rtype_string = "LA_CF";
      default : entries_0_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : entries_0_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_0_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_0_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_0_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : entries_0_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : entries_0_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_0_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_0_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_0_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : entries_0_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_immUsage)
      ImmUsageType_NONE : entries_0_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entries_0_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entries_0_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entries_0_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entries_0_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entries_0_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entries_0_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : entries_0_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : entries_0_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entries_0_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entries_0_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entries_0_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : entries_0_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_memCtrl_size)
      MemAccessSize_B : entries_0_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : entries_0_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : entries_0_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : entries_0_uop_decoded_memCtrl_size_string = "D";
      default : entries_0_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : entries_0_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entries_0_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entries_0_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entries_0_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entries_0_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entries_0_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entries_0_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entries_0_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entries_0_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entries_0_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entries_0_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entries_0_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entries_0_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entries_0_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entries_0_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entries_0_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entries_0_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entries_0_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entries_0_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entries_0_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entries_0_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entries_0_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_0_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_0_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_0_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entries_0_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : entries_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : entries_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : entries_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : entries_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : entries_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : entries_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : entries_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : entries_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : entries_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : entries_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : entries_0_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : entries_0_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : entries_0_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : entries_0_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : entries_0_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_0_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : entries_0_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : entries_0_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : entries_0_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : entries_0_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : entries_0_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_uopCode)
      BaseUopCode_NOP : entries_1_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : entries_1_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : entries_1_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : entries_1_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : entries_1_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : entries_1_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : entries_1_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : entries_1_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : entries_1_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : entries_1_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : entries_1_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : entries_1_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : entries_1_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : entries_1_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : entries_1_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : entries_1_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : entries_1_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : entries_1_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : entries_1_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : entries_1_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : entries_1_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : entries_1_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : entries_1_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : entries_1_uop_decoded_uopCode_string = "IDLE       ";
      default : entries_1_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_exeUnit)
      ExeUnitType_NONE : entries_1_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : entries_1_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : entries_1_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : entries_1_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : entries_1_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : entries_1_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : entries_1_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : entries_1_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : entries_1_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : entries_1_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_isa)
      IsaType_UNKNOWN : entries_1_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : entries_1_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : entries_1_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : entries_1_uop_decoded_isa_string = "LOONGARCH";
      default : entries_1_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_archDest_rtype)
      ArchRegType_GPR : entries_1_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_1_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_1_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_1_uop_decoded_archDest_rtype_string = "LA_CF";
      default : entries_1_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : entries_1_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_1_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_1_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_1_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : entries_1_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : entries_1_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_1_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_1_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_1_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : entries_1_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_immUsage)
      ImmUsageType_NONE : entries_1_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entries_1_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entries_1_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entries_1_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entries_1_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entries_1_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entries_1_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : entries_1_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : entries_1_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entries_1_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entries_1_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entries_1_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : entries_1_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_memCtrl_size)
      MemAccessSize_B : entries_1_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : entries_1_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : entries_1_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : entries_1_uop_decoded_memCtrl_size_string = "D";
      default : entries_1_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : entries_1_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entries_1_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entries_1_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entries_1_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entries_1_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entries_1_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entries_1_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entries_1_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entries_1_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entries_1_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entries_1_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entries_1_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entries_1_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entries_1_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entries_1_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entries_1_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entries_1_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entries_1_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entries_1_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entries_1_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entries_1_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entries_1_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_1_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_1_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_1_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entries_1_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : entries_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : entries_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : entries_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : entries_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : entries_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : entries_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : entries_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : entries_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : entries_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : entries_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : entries_1_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : entries_1_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : entries_1_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : entries_1_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : entries_1_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_1_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : entries_1_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : entries_1_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : entries_1_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : entries_1_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : entries_1_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_uopCode)
      BaseUopCode_NOP : entries_2_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : entries_2_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : entries_2_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : entries_2_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : entries_2_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : entries_2_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : entries_2_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : entries_2_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : entries_2_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : entries_2_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : entries_2_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : entries_2_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : entries_2_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : entries_2_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : entries_2_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : entries_2_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : entries_2_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : entries_2_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : entries_2_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : entries_2_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : entries_2_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : entries_2_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : entries_2_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : entries_2_uop_decoded_uopCode_string = "IDLE       ";
      default : entries_2_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_exeUnit)
      ExeUnitType_NONE : entries_2_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : entries_2_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : entries_2_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : entries_2_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : entries_2_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : entries_2_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : entries_2_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : entries_2_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : entries_2_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : entries_2_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_isa)
      IsaType_UNKNOWN : entries_2_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : entries_2_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : entries_2_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : entries_2_uop_decoded_isa_string = "LOONGARCH";
      default : entries_2_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_archDest_rtype)
      ArchRegType_GPR : entries_2_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_2_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_2_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_2_uop_decoded_archDest_rtype_string = "LA_CF";
      default : entries_2_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : entries_2_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_2_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_2_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_2_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : entries_2_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : entries_2_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_2_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_2_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_2_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : entries_2_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_immUsage)
      ImmUsageType_NONE : entries_2_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entries_2_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entries_2_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entries_2_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entries_2_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entries_2_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entries_2_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : entries_2_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : entries_2_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entries_2_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entries_2_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entries_2_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : entries_2_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_memCtrl_size)
      MemAccessSize_B : entries_2_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : entries_2_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : entries_2_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : entries_2_uop_decoded_memCtrl_size_string = "D";
      default : entries_2_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : entries_2_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entries_2_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entries_2_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entries_2_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entries_2_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entries_2_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entries_2_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entries_2_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entries_2_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entries_2_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entries_2_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entries_2_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entries_2_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entries_2_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entries_2_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entries_2_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entries_2_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entries_2_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entries_2_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entries_2_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entries_2_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entries_2_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_2_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_2_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_2_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entries_2_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : entries_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : entries_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : entries_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : entries_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : entries_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : entries_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : entries_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : entries_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : entries_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : entries_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : entries_2_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : entries_2_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : entries_2_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : entries_2_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : entries_2_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_2_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : entries_2_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : entries_2_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : entries_2_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : entries_2_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : entries_2_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_uopCode)
      BaseUopCode_NOP : entries_3_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : entries_3_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : entries_3_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : entries_3_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : entries_3_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : entries_3_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : entries_3_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : entries_3_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : entries_3_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : entries_3_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : entries_3_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : entries_3_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : entries_3_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : entries_3_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : entries_3_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : entries_3_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : entries_3_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : entries_3_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : entries_3_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : entries_3_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : entries_3_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : entries_3_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : entries_3_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : entries_3_uop_decoded_uopCode_string = "IDLE       ";
      default : entries_3_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_exeUnit)
      ExeUnitType_NONE : entries_3_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : entries_3_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : entries_3_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : entries_3_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : entries_3_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : entries_3_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : entries_3_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : entries_3_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : entries_3_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : entries_3_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_isa)
      IsaType_UNKNOWN : entries_3_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : entries_3_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : entries_3_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : entries_3_uop_decoded_isa_string = "LOONGARCH";
      default : entries_3_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_archDest_rtype)
      ArchRegType_GPR : entries_3_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_3_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_3_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_3_uop_decoded_archDest_rtype_string = "LA_CF";
      default : entries_3_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : entries_3_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_3_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_3_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_3_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : entries_3_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : entries_3_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_3_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_3_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_3_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : entries_3_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_immUsage)
      ImmUsageType_NONE : entries_3_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entries_3_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entries_3_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entries_3_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entries_3_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entries_3_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entries_3_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : entries_3_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : entries_3_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entries_3_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entries_3_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entries_3_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : entries_3_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_memCtrl_size)
      MemAccessSize_B : entries_3_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : entries_3_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : entries_3_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : entries_3_uop_decoded_memCtrl_size_string = "D";
      default : entries_3_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : entries_3_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entries_3_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entries_3_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entries_3_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entries_3_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entries_3_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entries_3_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entries_3_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entries_3_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entries_3_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entries_3_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entries_3_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entries_3_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entries_3_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entries_3_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entries_3_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entries_3_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entries_3_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entries_3_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entries_3_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entries_3_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entries_3_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entries_3_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entries_3_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entries_3_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entries_3_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : entries_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : entries_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : entries_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : entries_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : entries_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : entries_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : entries_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : entries_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : entries_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : entries_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : entries_3_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : entries_3_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : entries_3_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : entries_3_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : entries_3_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(entries_3_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : entries_3_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : entries_3_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : entries_3_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : entries_3_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : entries_3_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : _zz_io_issueOut_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : _zz_io_issueOut_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_isa)
      IsaType_UNKNOWN : _zz_io_issueOut_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : _zz_io_issueOut_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : _zz_io_issueOut_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : _zz_io_issueOut_payload_uop_decoded_isa_string = "LOONGARCH";
      default : _zz_io_issueOut_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : _zz_io_issueOut_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_issueOut_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_issueOut_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_issueOut_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : _zz_io_issueOut_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : _zz_io_issueOut_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_io_issueOut_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_io_issueOut_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_io_issueOut_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_io_issueOut_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_io_issueOut_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_io_issueOut_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : _zz_io_issueOut_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : _zz_io_issueOut_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : _zz_io_issueOut_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : _zz_io_issueOut_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : _zz_io_issueOut_payload_uop_decoded_memCtrl_size_string = "D";
      default : _zz_io_issueOut_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_uopCode)
      BaseUopCode_NOP : entriesNext_0_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : entriesNext_0_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : entriesNext_0_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : entriesNext_0_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : entriesNext_0_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : entriesNext_0_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : entriesNext_0_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : entriesNext_0_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : entriesNext_0_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : entriesNext_0_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : entriesNext_0_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : entriesNext_0_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : entriesNext_0_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : entriesNext_0_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : entriesNext_0_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : entriesNext_0_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : entriesNext_0_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : entriesNext_0_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : entriesNext_0_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : entriesNext_0_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : entriesNext_0_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : entriesNext_0_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : entriesNext_0_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : entriesNext_0_uop_decoded_uopCode_string = "IDLE       ";
      default : entriesNext_0_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_exeUnit)
      ExeUnitType_NONE : entriesNext_0_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : entriesNext_0_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : entriesNext_0_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : entriesNext_0_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : entriesNext_0_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : entriesNext_0_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : entriesNext_0_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : entriesNext_0_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : entriesNext_0_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : entriesNext_0_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_isa)
      IsaType_UNKNOWN : entriesNext_0_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : entriesNext_0_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : entriesNext_0_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : entriesNext_0_uop_decoded_isa_string = "LOONGARCH";
      default : entriesNext_0_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_archDest_rtype)
      ArchRegType_GPR : entriesNext_0_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_0_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_0_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_0_uop_decoded_archDest_rtype_string = "LA_CF";
      default : entriesNext_0_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : entriesNext_0_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_0_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_0_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_0_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : entriesNext_0_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : entriesNext_0_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_0_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_0_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_0_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : entriesNext_0_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_immUsage)
      ImmUsageType_NONE : entriesNext_0_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entriesNext_0_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entriesNext_0_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entriesNext_0_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entriesNext_0_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entriesNext_0_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entriesNext_0_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : entriesNext_0_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : entriesNext_0_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entriesNext_0_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entriesNext_0_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entriesNext_0_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : entriesNext_0_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_memCtrl_size)
      MemAccessSize_B : entriesNext_0_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : entriesNext_0_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : entriesNext_0_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : entriesNext_0_uop_decoded_memCtrl_size_string = "D";
      default : entriesNext_0_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : entriesNext_0_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entriesNext_0_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entriesNext_0_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entriesNext_0_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entriesNext_0_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entriesNext_0_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entriesNext_0_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entriesNext_0_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entriesNext_0_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entriesNext_0_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entriesNext_0_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entriesNext_0_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entriesNext_0_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entriesNext_0_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entriesNext_0_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entriesNext_0_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entriesNext_0_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entriesNext_0_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entriesNext_0_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entriesNext_0_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entriesNext_0_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : entriesNext_0_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : entriesNext_0_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : entriesNext_0_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : entriesNext_0_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : entriesNext_0_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_uopCode)
      BaseUopCode_NOP : entriesNext_1_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : entriesNext_1_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : entriesNext_1_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : entriesNext_1_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : entriesNext_1_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : entriesNext_1_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : entriesNext_1_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : entriesNext_1_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : entriesNext_1_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : entriesNext_1_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : entriesNext_1_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : entriesNext_1_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : entriesNext_1_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : entriesNext_1_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : entriesNext_1_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : entriesNext_1_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : entriesNext_1_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : entriesNext_1_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : entriesNext_1_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : entriesNext_1_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : entriesNext_1_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : entriesNext_1_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : entriesNext_1_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : entriesNext_1_uop_decoded_uopCode_string = "IDLE       ";
      default : entriesNext_1_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_exeUnit)
      ExeUnitType_NONE : entriesNext_1_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : entriesNext_1_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : entriesNext_1_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : entriesNext_1_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : entriesNext_1_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : entriesNext_1_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : entriesNext_1_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : entriesNext_1_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : entriesNext_1_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : entriesNext_1_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_isa)
      IsaType_UNKNOWN : entriesNext_1_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : entriesNext_1_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : entriesNext_1_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : entriesNext_1_uop_decoded_isa_string = "LOONGARCH";
      default : entriesNext_1_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_archDest_rtype)
      ArchRegType_GPR : entriesNext_1_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_1_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_1_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_1_uop_decoded_archDest_rtype_string = "LA_CF";
      default : entriesNext_1_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : entriesNext_1_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_1_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_1_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_1_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : entriesNext_1_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : entriesNext_1_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_1_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_1_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_1_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : entriesNext_1_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_immUsage)
      ImmUsageType_NONE : entriesNext_1_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entriesNext_1_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entriesNext_1_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entriesNext_1_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entriesNext_1_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entriesNext_1_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entriesNext_1_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : entriesNext_1_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : entriesNext_1_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entriesNext_1_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entriesNext_1_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entriesNext_1_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : entriesNext_1_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_memCtrl_size)
      MemAccessSize_B : entriesNext_1_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : entriesNext_1_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : entriesNext_1_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : entriesNext_1_uop_decoded_memCtrl_size_string = "D";
      default : entriesNext_1_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : entriesNext_1_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entriesNext_1_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entriesNext_1_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entriesNext_1_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entriesNext_1_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entriesNext_1_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entriesNext_1_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entriesNext_1_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entriesNext_1_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entriesNext_1_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entriesNext_1_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entriesNext_1_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entriesNext_1_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entriesNext_1_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entriesNext_1_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entriesNext_1_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entriesNext_1_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entriesNext_1_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entriesNext_1_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entriesNext_1_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entriesNext_1_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : entriesNext_1_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : entriesNext_1_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : entriesNext_1_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : entriesNext_1_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : entriesNext_1_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_uopCode)
      BaseUopCode_NOP : entriesNext_2_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : entriesNext_2_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : entriesNext_2_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : entriesNext_2_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : entriesNext_2_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : entriesNext_2_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : entriesNext_2_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : entriesNext_2_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : entriesNext_2_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : entriesNext_2_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : entriesNext_2_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : entriesNext_2_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : entriesNext_2_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : entriesNext_2_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : entriesNext_2_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : entriesNext_2_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : entriesNext_2_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : entriesNext_2_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : entriesNext_2_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : entriesNext_2_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : entriesNext_2_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : entriesNext_2_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : entriesNext_2_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : entriesNext_2_uop_decoded_uopCode_string = "IDLE       ";
      default : entriesNext_2_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_exeUnit)
      ExeUnitType_NONE : entriesNext_2_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : entriesNext_2_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : entriesNext_2_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : entriesNext_2_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : entriesNext_2_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : entriesNext_2_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : entriesNext_2_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : entriesNext_2_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : entriesNext_2_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : entriesNext_2_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_isa)
      IsaType_UNKNOWN : entriesNext_2_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : entriesNext_2_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : entriesNext_2_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : entriesNext_2_uop_decoded_isa_string = "LOONGARCH";
      default : entriesNext_2_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_archDest_rtype)
      ArchRegType_GPR : entriesNext_2_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_2_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_2_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_2_uop_decoded_archDest_rtype_string = "LA_CF";
      default : entriesNext_2_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : entriesNext_2_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_2_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_2_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_2_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : entriesNext_2_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : entriesNext_2_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_2_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_2_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_2_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : entriesNext_2_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_immUsage)
      ImmUsageType_NONE : entriesNext_2_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entriesNext_2_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entriesNext_2_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entriesNext_2_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entriesNext_2_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entriesNext_2_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entriesNext_2_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : entriesNext_2_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : entriesNext_2_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entriesNext_2_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entriesNext_2_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entriesNext_2_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : entriesNext_2_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_memCtrl_size)
      MemAccessSize_B : entriesNext_2_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : entriesNext_2_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : entriesNext_2_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : entriesNext_2_uop_decoded_memCtrl_size_string = "D";
      default : entriesNext_2_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : entriesNext_2_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entriesNext_2_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entriesNext_2_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entriesNext_2_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entriesNext_2_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entriesNext_2_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entriesNext_2_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entriesNext_2_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entriesNext_2_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entriesNext_2_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entriesNext_2_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entriesNext_2_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entriesNext_2_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entriesNext_2_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entriesNext_2_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entriesNext_2_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entriesNext_2_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entriesNext_2_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entriesNext_2_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entriesNext_2_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entriesNext_2_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : entriesNext_2_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : entriesNext_2_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : entriesNext_2_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : entriesNext_2_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : entriesNext_2_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_uopCode)
      BaseUopCode_NOP : entriesNext_3_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : entriesNext_3_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : entriesNext_3_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : entriesNext_3_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : entriesNext_3_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : entriesNext_3_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : entriesNext_3_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : entriesNext_3_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : entriesNext_3_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : entriesNext_3_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : entriesNext_3_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : entriesNext_3_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : entriesNext_3_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : entriesNext_3_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : entriesNext_3_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : entriesNext_3_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : entriesNext_3_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : entriesNext_3_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : entriesNext_3_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : entriesNext_3_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : entriesNext_3_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : entriesNext_3_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : entriesNext_3_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : entriesNext_3_uop_decoded_uopCode_string = "IDLE       ";
      default : entriesNext_3_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_exeUnit)
      ExeUnitType_NONE : entriesNext_3_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : entriesNext_3_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : entriesNext_3_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : entriesNext_3_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : entriesNext_3_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : entriesNext_3_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : entriesNext_3_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : entriesNext_3_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : entriesNext_3_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : entriesNext_3_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_isa)
      IsaType_UNKNOWN : entriesNext_3_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : entriesNext_3_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : entriesNext_3_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : entriesNext_3_uop_decoded_isa_string = "LOONGARCH";
      default : entriesNext_3_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_archDest_rtype)
      ArchRegType_GPR : entriesNext_3_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_3_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_3_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_3_uop_decoded_archDest_rtype_string = "LA_CF";
      default : entriesNext_3_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : entriesNext_3_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_3_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_3_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_3_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : entriesNext_3_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : entriesNext_3_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_3_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_3_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_3_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : entriesNext_3_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_immUsage)
      ImmUsageType_NONE : entriesNext_3_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entriesNext_3_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entriesNext_3_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entriesNext_3_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entriesNext_3_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entriesNext_3_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entriesNext_3_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : entriesNext_3_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : entriesNext_3_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entriesNext_3_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entriesNext_3_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entriesNext_3_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : entriesNext_3_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_memCtrl_size)
      MemAccessSize_B : entriesNext_3_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : entriesNext_3_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : entriesNext_3_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : entriesNext_3_uop_decoded_memCtrl_size_string = "D";
      default : entriesNext_3_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : entriesNext_3_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : entriesNext_3_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : entriesNext_3_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : entriesNext_3_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : entriesNext_3_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : entriesNext_3_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : entriesNext_3_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : entriesNext_3_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : entriesNext_3_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : entriesNext_3_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : entriesNext_3_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : entriesNext_3_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : entriesNext_3_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : entriesNext_3_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : entriesNext_3_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : entriesNext_3_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : entriesNext_3_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : entriesNext_3_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : entriesNext_3_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : entriesNext_3_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : entriesNext_3_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : entriesNext_3_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : entriesNext_3_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : entriesNext_3_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : entriesNext_3_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : entriesNext_3_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  `endif

  assign io_issueOut_fire = (io_issueOut_valid && io_issueOut_ready);
  assign localWakeupValid = (io_issueOut_fire && io_issueOut_payload_writesToPhysReg);
  always @(*) begin
    wokeUpSrc1Mask = 4'b0000;
    if(entryValids_0) begin
      if(when_IssueQueueComponent_l103) begin
        wokeUpSrc1Mask[0] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_1) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_2) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_3) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_4) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
    end
    if(entryValids_1) begin
      if(when_IssueQueueComponent_l103_1) begin
        wokeUpSrc1Mask[1] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_5) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_6) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_7) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_8) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_9) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
    end
    if(entryValids_2) begin
      if(when_IssueQueueComponent_l103_2) begin
        wokeUpSrc1Mask[2] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_10) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_11) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_12) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_13) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_14) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
    end
    if(entryValids_3) begin
      if(when_IssueQueueComponent_l103_3) begin
        wokeUpSrc1Mask[3] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_15) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_16) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_17) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_18) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_19) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    wokeUpSrc2Mask = 4'b0000;
    if(entryValids_0) begin
      if(when_IssueQueueComponent_l106) begin
        wokeUpSrc2Mask[0] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_1) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_2) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_3) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_4) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
    end
    if(entryValids_1) begin
      if(when_IssueQueueComponent_l106_1) begin
        wokeUpSrc2Mask[1] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_5) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_6) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_7) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_8) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_9) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
    end
    if(entryValids_2) begin
      if(when_IssueQueueComponent_l106_2) begin
        wokeUpSrc2Mask[2] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_10) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_11) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_12) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_13) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_14) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
    end
    if(entryValids_3) begin
      if(when_IssueQueueComponent_l106_3) begin
        wokeUpSrc2Mask[3] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_15) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_16) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_17) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_18) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_19) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
    end
  end

  assign _zz_when_IssueQueueComponent_l103 = ((! entries_0_src1Ready) && entries_0_useSrc1);
  assign _zz_when_IssueQueueComponent_l106 = ((! entries_0_src2Ready) && entries_0_useSrc2);
  assign when_IssueQueueComponent_l103 = ((_zz_when_IssueQueueComponent_l103 && localWakeupValid) && (entries_0_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106 = ((_zz_when_IssueQueueComponent_l106 && localWakeupValid) && (entries_0_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_1 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_1 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_2 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_2 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_3 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_3 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_4 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_4 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_1 = ((! entries_1_src1Ready) && entries_1_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_1 = ((! entries_1_src2Ready) && entries_1_useSrc2);
  assign when_IssueQueueComponent_l103_1 = ((_zz_when_IssueQueueComponent_l103_1 && localWakeupValid) && (entries_1_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_1 = ((_zz_when_IssueQueueComponent_l106_1 && localWakeupValid) && (entries_1_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_5 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_5 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_6 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_6 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_7 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_7 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_8 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_8 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_9 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_9 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_2 = ((! entries_2_src1Ready) && entries_2_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_2 = ((! entries_2_src2Ready) && entries_2_useSrc2);
  assign when_IssueQueueComponent_l103_2 = ((_zz_when_IssueQueueComponent_l103_2 && localWakeupValid) && (entries_2_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_2 = ((_zz_when_IssueQueueComponent_l106_2 && localWakeupValid) && (entries_2_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_10 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_10 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_11 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_11 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_12 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_12 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_13 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_13 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_14 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_14 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_3 = ((! entries_3_src1Ready) && entries_3_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_3 = ((! entries_3_src2Ready) && entries_3_useSrc2);
  assign when_IssueQueueComponent_l103_3 = ((_zz_when_IssueQueueComponent_l103_3 && localWakeupValid) && (entries_3_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_3 = ((_zz_when_IssueQueueComponent_l106_3 && localWakeupValid) && (entries_3_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_15 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_15 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_16 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_16 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_17 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_17 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_18 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_18 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_19 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_19 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign entriesReadyToIssue_0 = ((entryValids_0 && ((! entries_0_useSrc1) || entries_0_src1Ready)) && ((! entries_0_useSrc2) || entries_0_src2Ready));
  assign entriesReadyToIssue_1 = ((entryValids_1 && ((! entries_1_useSrc1) || entries_1_src1Ready)) && ((! entries_1_useSrc2) || entries_1_src2Ready));
  assign entriesReadyToIssue_2 = ((entryValids_2 && ((! entries_2_useSrc1) || entries_2_src1Ready)) && ((! entries_2_useSrc2) || entries_2_src2Ready));
  assign entriesReadyToIssue_3 = ((entryValids_3 && ((! entries_3_useSrc1) || entries_3_src1Ready)) && ((! entries_3_useSrc2) || entries_3_src2Ready));
  assign issueRequestMask = {entriesReadyToIssue_3,{entriesReadyToIssue_2,{entriesReadyToIssue_1,entriesReadyToIssue_0}}};
  assign issueRequestMask_ohFirst_input = issueRequestMask;
  assign issueRequestMask_ohFirst_masked = (issueRequestMask_ohFirst_input & (~ _zz_issueRequestMask_ohFirst_masked));
  assign issueRequestOh = issueRequestMask_ohFirst_masked;
  assign _zz_issueIdx = issueRequestOh[3];
  assign _zz_issueIdx_1 = (issueRequestOh[1] || _zz_issueIdx);
  assign _zz_issueIdx_2 = (issueRequestOh[2] || _zz_issueIdx);
  assign issueIdx = {_zz_issueIdx_2,_zz_issueIdx_1};
  assign io_issueOut_valid = ((|issueRequestOh) && (! io_flush));
  assign _zz_io_issueOut_payload_uop_decoded_uopCode = _zz__zz_io_issueOut_payload_uop_decoded_uopCode;
  assign _zz_io_issueOut_payload_uop_decoded_exeUnit = _zz__zz_io_issueOut_payload_uop_decoded_exeUnit;
  assign _zz_io_issueOut_payload_uop_decoded_isa = _zz__zz_io_issueOut_payload_uop_decoded_isa;
  assign _zz_io_issueOut_payload_uop_decoded_archDest_rtype = _zz__zz_io_issueOut_payload_uop_decoded_archDest_rtype;
  assign _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype = _zz__zz_io_issueOut_payload_uop_decoded_archSrc1_rtype;
  assign _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype = _zz__zz_io_issueOut_payload_uop_decoded_archSrc2_rtype;
  assign _zz_io_issueOut_payload_uop_decoded_immUsage = _zz__zz_io_issueOut_payload_uop_decoded_immUsage;
  assign _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp = _zz__zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp;
  assign _zz_io_issueOut_payload_uop_decoded_memCtrl_size = _zz__zz_io_issueOut_payload_uop_decoded_memCtrl_size;
  assign _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition = _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_condition;
  assign _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype = _zz__zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype;
  assign _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  assign _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  assign _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest = _zz__zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest;
  assign _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode = _zz__zz_io_issueOut_payload_uop_decoded_decodeExceptionCode;
  assign io_issueOut_payload_uop_decoded_pc = _zz_io_issueOut_payload_uop_decoded_pc;
  assign io_issueOut_payload_uop_decoded_isValid = _zz_io_issueOut_payload_uop_decoded_isValid;
  assign io_issueOut_payload_uop_decoded_uopCode = _zz_io_issueOut_payload_uop_decoded_uopCode;
  assign io_issueOut_payload_uop_decoded_exeUnit = _zz_io_issueOut_payload_uop_decoded_exeUnit;
  assign io_issueOut_payload_uop_decoded_isa = _zz_io_issueOut_payload_uop_decoded_isa;
  assign io_issueOut_payload_uop_decoded_archDest_idx = _zz_io_issueOut_payload_uop_decoded_archDest_idx;
  assign io_issueOut_payload_uop_decoded_archDest_rtype = _zz_io_issueOut_payload_uop_decoded_archDest_rtype;
  assign io_issueOut_payload_uop_decoded_writeArchDestEn = _zz_io_issueOut_payload_uop_decoded_writeArchDestEn;
  assign io_issueOut_payload_uop_decoded_archSrc1_idx = _zz_io_issueOut_payload_uop_decoded_archSrc1_idx;
  assign io_issueOut_payload_uop_decoded_archSrc1_rtype = _zz_io_issueOut_payload_uop_decoded_archSrc1_rtype;
  assign io_issueOut_payload_uop_decoded_useArchSrc1 = _zz_io_issueOut_payload_uop_decoded_useArchSrc1;
  assign io_issueOut_payload_uop_decoded_archSrc2_idx = _zz_io_issueOut_payload_uop_decoded_archSrc2_idx;
  assign io_issueOut_payload_uop_decoded_archSrc2_rtype = _zz_io_issueOut_payload_uop_decoded_archSrc2_rtype;
  assign io_issueOut_payload_uop_decoded_useArchSrc2 = _zz_io_issueOut_payload_uop_decoded_useArchSrc2;
  assign io_issueOut_payload_uop_decoded_usePcForAddr = _zz_io_issueOut_payload_uop_decoded_usePcForAddr;
  assign io_issueOut_payload_uop_decoded_imm = _zz_io_issueOut_payload_uop_decoded_imm;
  assign io_issueOut_payload_uop_decoded_immUsage = _zz_io_issueOut_payload_uop_decoded_immUsage;
  assign io_issueOut_payload_uop_decoded_aluCtrl_valid = _zz_io_issueOut_payload_uop_decoded_aluCtrl_valid;
  assign io_issueOut_payload_uop_decoded_aluCtrl_isSub = _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSub;
  assign io_issueOut_payload_uop_decoded_aluCtrl_isAdd = _zz_io_issueOut_payload_uop_decoded_aluCtrl_isAdd;
  assign io_issueOut_payload_uop_decoded_aluCtrl_isSigned = _zz_io_issueOut_payload_uop_decoded_aluCtrl_isSigned;
  assign io_issueOut_payload_uop_decoded_aluCtrl_logicOp = _zz_io_issueOut_payload_uop_decoded_aluCtrl_logicOp;
  assign io_issueOut_payload_uop_decoded_shiftCtrl_valid = _zz_io_issueOut_payload_uop_decoded_shiftCtrl_valid;
  assign io_issueOut_payload_uop_decoded_shiftCtrl_isRight = _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRight;
  assign io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic = _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isArithmetic;
  assign io_issueOut_payload_uop_decoded_shiftCtrl_isRotate = _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isRotate;
  assign io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord = _zz_io_issueOut_payload_uop_decoded_shiftCtrl_isDoubleWord;
  assign io_issueOut_payload_uop_decoded_mulDivCtrl_valid = _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_valid;
  assign io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv = _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isDiv;
  assign io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned = _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isSigned;
  assign io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp = _zz_io_issueOut_payload_uop_decoded_mulDivCtrl_isWordOp;
  assign io_issueOut_payload_uop_decoded_memCtrl_size = _zz_io_issueOut_payload_uop_decoded_memCtrl_size;
  assign io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad = _zz_io_issueOut_payload_uop_decoded_memCtrl_isSignedLoad;
  assign io_issueOut_payload_uop_decoded_memCtrl_isStore = _zz_io_issueOut_payload_uop_decoded_memCtrl_isStore;
  assign io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked = _zz_io_issueOut_payload_uop_decoded_memCtrl_isLoadLinked;
  assign io_issueOut_payload_uop_decoded_memCtrl_isStoreCond = _zz_io_issueOut_payload_uop_decoded_memCtrl_isStoreCond;
  assign io_issueOut_payload_uop_decoded_memCtrl_atomicOp = _zz_io_issueOut_payload_uop_decoded_memCtrl_atomicOp;
  assign io_issueOut_payload_uop_decoded_memCtrl_isFence = _zz_io_issueOut_payload_uop_decoded_memCtrl_isFence;
  assign io_issueOut_payload_uop_decoded_memCtrl_fenceMode = _zz_io_issueOut_payload_uop_decoded_memCtrl_fenceMode;
  assign io_issueOut_payload_uop_decoded_memCtrl_isCacheOp = _zz_io_issueOut_payload_uop_decoded_memCtrl_isCacheOp;
  assign io_issueOut_payload_uop_decoded_memCtrl_cacheOpType = _zz_io_issueOut_payload_uop_decoded_memCtrl_cacheOpType;
  assign io_issueOut_payload_uop_decoded_memCtrl_isPrefetch = _zz_io_issueOut_payload_uop_decoded_memCtrl_isPrefetch;
  assign io_issueOut_payload_uop_decoded_branchCtrl_condition = _zz_io_issueOut_payload_uop_decoded_branchCtrl_condition;
  assign io_issueOut_payload_uop_decoded_branchCtrl_isJump = _zz_io_issueOut_payload_uop_decoded_branchCtrl_isJump;
  assign io_issueOut_payload_uop_decoded_branchCtrl_isLink = _zz_io_issueOut_payload_uop_decoded_branchCtrl_isLink;
  assign io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx = _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_idx;
  assign io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype = _zz_io_issueOut_payload_uop_decoded_branchCtrl_linkReg_rtype;
  assign io_issueOut_payload_uop_decoded_branchCtrl_isIndirect = _zz_io_issueOut_payload_uop_decoded_branchCtrl_isIndirect;
  assign io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx = _zz_io_issueOut_payload_uop_decoded_branchCtrl_laCfIdx;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_opType = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_opType;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fpSizeDest;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_roundingMode;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isIntegerDest;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_isSignedCvt;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
  assign io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond = _zz_io_issueOut_payload_uop_decoded_fpuCtrl_fcmpCond;
  assign io_issueOut_payload_uop_decoded_csrCtrl_csrAddr = _zz_io_issueOut_payload_uop_decoded_csrCtrl_csrAddr;
  assign io_issueOut_payload_uop_decoded_csrCtrl_isWrite = _zz_io_issueOut_payload_uop_decoded_csrCtrl_isWrite;
  assign io_issueOut_payload_uop_decoded_csrCtrl_isRead = _zz_io_issueOut_payload_uop_decoded_csrCtrl_isRead;
  assign io_issueOut_payload_uop_decoded_csrCtrl_isExchange = _zz_io_issueOut_payload_uop_decoded_csrCtrl_isExchange;
  assign io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc = _zz_io_issueOut_payload_uop_decoded_csrCtrl_useUimmAsSrc;
  assign io_issueOut_payload_uop_decoded_sysCtrl_sysCode = _zz_io_issueOut_payload_uop_decoded_sysCtrl_sysCode;
  assign io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn = _zz_io_issueOut_payload_uop_decoded_sysCtrl_isExceptionReturn;
  assign io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp = _zz_io_issueOut_payload_uop_decoded_sysCtrl_isTlbOp;
  assign io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType = _zz_io_issueOut_payload_uop_decoded_sysCtrl_tlbOpType;
  assign io_issueOut_payload_uop_decoded_decodeExceptionCode = _zz_io_issueOut_payload_uop_decoded_decodeExceptionCode;
  assign io_issueOut_payload_uop_decoded_hasDecodeException = _zz_io_issueOut_payload_uop_decoded_hasDecodeException;
  assign io_issueOut_payload_uop_decoded_isMicrocode = _zz_io_issueOut_payload_uop_decoded_isMicrocode;
  assign io_issueOut_payload_uop_decoded_microcodeEntry = _zz_io_issueOut_payload_uop_decoded_microcodeEntry;
  assign io_issueOut_payload_uop_decoded_isSerializing = _zz_io_issueOut_payload_uop_decoded_isSerializing;
  assign io_issueOut_payload_uop_decoded_isBranchOrJump = _zz_io_issueOut_payload_uop_decoded_isBranchOrJump;
  assign io_issueOut_payload_uop_decoded_branchPrediction_isTaken = _zz_io_issueOut_payload_uop_decoded_branchPrediction_isTaken;
  assign io_issueOut_payload_uop_decoded_branchPrediction_target = _zz_io_issueOut_payload_uop_decoded_branchPrediction_target;
  assign io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted = _zz_io_issueOut_payload_uop_decoded_branchPrediction_wasPredicted;
  assign io_issueOut_payload_uop_rename_physSrc1_idx = _zz_io_issueOut_payload_uop_rename_physSrc1_idx;
  assign io_issueOut_payload_uop_rename_physSrc1IsFpr = _zz_io_issueOut_payload_uop_rename_physSrc1IsFpr;
  assign io_issueOut_payload_uop_rename_physSrc2_idx = _zz_io_issueOut_payload_uop_rename_physSrc2_idx;
  assign io_issueOut_payload_uop_rename_physSrc2IsFpr = _zz_io_issueOut_payload_uop_rename_physSrc2IsFpr;
  assign io_issueOut_payload_uop_rename_physDest_idx = _zz_io_issueOut_payload_uop_rename_physDest_idx;
  assign io_issueOut_payload_uop_rename_physDestIsFpr = _zz_io_issueOut_payload_uop_rename_physDestIsFpr;
  assign io_issueOut_payload_uop_rename_oldPhysDest_idx = _zz_io_issueOut_payload_uop_rename_oldPhysDest_idx;
  assign io_issueOut_payload_uop_rename_oldPhysDestIsFpr = _zz_io_issueOut_payload_uop_rename_oldPhysDestIsFpr;
  assign io_issueOut_payload_uop_rename_allocatesPhysDest = _zz_io_issueOut_payload_uop_rename_allocatesPhysDest;
  assign io_issueOut_payload_uop_rename_writesToPhysReg = _zz_io_issueOut_payload_uop_rename_writesToPhysReg;
  assign io_issueOut_payload_uop_robPtr = _zz_io_issueOut_payload_uop_robPtr;
  assign io_issueOut_payload_uop_uniqueId = _zz_io_issueOut_payload_uop_uniqueId;
  assign io_issueOut_payload_uop_dispatched = _zz_io_issueOut_payload_uop_dispatched;
  assign io_issueOut_payload_uop_executed = _zz_io_issueOut_payload_uop_executed;
  assign io_issueOut_payload_uop_hasException = _zz_io_issueOut_payload_uop_hasException;
  assign io_issueOut_payload_uop_exceptionCode = _zz_io_issueOut_payload_uop_exceptionCode;
  assign io_issueOut_payload_robPtr = _zz_io_issueOut_payload_robPtr;
  assign io_issueOut_payload_physDest_idx = _zz_io_issueOut_payload_physDest_idx;
  assign io_issueOut_payload_physDestIsFpr = _zz_io_issueOut_payload_physDestIsFpr;
  assign io_issueOut_payload_writesToPhysReg = _zz_io_issueOut_payload_writesToPhysReg;
  assign io_issueOut_payload_useSrc1 = _zz_io_issueOut_payload_useSrc1;
  assign io_issueOut_payload_src1Data = _zz_io_issueOut_payload_src1Data;
  assign io_issueOut_payload_src1Tag = _zz_io_issueOut_payload_src1Tag;
  assign io_issueOut_payload_src1Ready = _zz_io_issueOut_payload_src1Ready;
  assign io_issueOut_payload_src1IsFpr = _zz_io_issueOut_payload_src1IsFpr;
  assign io_issueOut_payload_useSrc2 = _zz_io_issueOut_payload_useSrc2;
  assign io_issueOut_payload_src2Data = _zz_io_issueOut_payload_src2Data;
  assign io_issueOut_payload_src2Tag = _zz_io_issueOut_payload_src2Tag;
  assign io_issueOut_payload_src2Ready = _zz_io_issueOut_payload_src2Ready;
  assign io_issueOut_payload_src2IsFpr = _zz_io_issueOut_payload_src2IsFpr;
  assign io_issueOut_payload_mulDivCtrl_valid = _zz_io_issueOut_payload_mulDivCtrl_valid;
  assign io_issueOut_payload_mulDivCtrl_isDiv = _zz_io_issueOut_payload_mulDivCtrl_isDiv;
  assign io_issueOut_payload_mulDivCtrl_isSigned = _zz_io_issueOut_payload_mulDivCtrl_isSigned;
  assign io_issueOut_payload_mulDivCtrl_isWordOp = _zz_io_issueOut_payload_mulDivCtrl_isWordOp;
  assign freeSlotsMask = {(! entryValids_3),{(! entryValids_2),{(! entryValids_1),(! entryValids_0)}}};
  assign hasSpaceForNewEntry = ((|freeSlotsMask) || io_issueOut_fire);
  assign io_allocateIn_ready = (hasSpaceForNewEntry && (! io_flush));
  always @(*) begin
    firedSlotMask = 4'b0000;
    if(io_issueOut_fire) begin
      firedSlotMask[issueIdx] = 1'b1;
    end
  end

  assign _zz_allocationMask = (freeSlotsMask | firedSlotMask);
  assign allocationMask = (_zz_allocationMask & (~ _zz_allocationMask_1));
  assign _zz_allocateIdx = allocationMask[3];
  assign _zz_allocateIdx_1 = (allocationMask[1] || _zz_allocateIdx);
  assign _zz_allocateIdx_2 = (allocationMask[2] || _zz_allocateIdx);
  assign allocateIdx = {_zz_allocateIdx_2,_zz_allocateIdx_1};
  always @(*) begin
    entriesNext_0_uop_decoded_pc = entries_0_uop_decoded_pc;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_pc = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_isValid = entries_0_uop_decoded_isValid;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_isValid = io_allocateIn_payload_uop_decoded_isValid;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_uopCode = entries_0_uop_decoded_uopCode;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_uopCode = io_allocateIn_payload_uop_decoded_uopCode;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_exeUnit = entries_0_uop_decoded_exeUnit;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_exeUnit = io_allocateIn_payload_uop_decoded_exeUnit;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_isa = entries_0_uop_decoded_isa;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_isa = io_allocateIn_payload_uop_decoded_isa;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_archDest_idx = entries_0_uop_decoded_archDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_archDest_idx = io_allocateIn_payload_uop_decoded_archDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_archDest_rtype = entries_0_uop_decoded_archDest_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_archDest_rtype = io_allocateIn_payload_uop_decoded_archDest_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_writeArchDestEn = entries_0_uop_decoded_writeArchDestEn;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_writeArchDestEn = io_allocateIn_payload_uop_decoded_writeArchDestEn;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_archSrc1_idx = entries_0_uop_decoded_archSrc1_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_archSrc1_idx = io_allocateIn_payload_uop_decoded_archSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_archSrc1_rtype = entries_0_uop_decoded_archSrc1_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_archSrc1_rtype = io_allocateIn_payload_uop_decoded_archSrc1_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_useArchSrc1 = entries_0_uop_decoded_useArchSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_useArchSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_archSrc2_idx = entries_0_uop_decoded_archSrc2_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_archSrc2_idx = io_allocateIn_payload_uop_decoded_archSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_archSrc2_rtype = entries_0_uop_decoded_archSrc2_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_archSrc2_rtype = io_allocateIn_payload_uop_decoded_archSrc2_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_useArchSrc2 = entries_0_uop_decoded_useArchSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_useArchSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_usePcForAddr = entries_0_uop_decoded_usePcForAddr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_usePcForAddr = io_allocateIn_payload_uop_decoded_usePcForAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_imm = entries_0_uop_decoded_imm;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_immUsage = entries_0_uop_decoded_immUsage;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_immUsage = io_allocateIn_payload_uop_decoded_immUsage;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_aluCtrl_valid = entries_0_uop_decoded_aluCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_aluCtrl_valid = io_allocateIn_payload_uop_decoded_aluCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_aluCtrl_isSub = entries_0_uop_decoded_aluCtrl_isSub;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_aluCtrl_isSub = io_allocateIn_payload_uop_decoded_aluCtrl_isSub;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_aluCtrl_isAdd = entries_0_uop_decoded_aluCtrl_isAdd;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_aluCtrl_isAdd = io_allocateIn_payload_uop_decoded_aluCtrl_isAdd;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_aluCtrl_isSigned = entries_0_uop_decoded_aluCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_aluCtrl_isSigned = io_allocateIn_payload_uop_decoded_aluCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_aluCtrl_logicOp = entries_0_uop_decoded_aluCtrl_logicOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_aluCtrl_logicOp = io_allocateIn_payload_uop_decoded_aluCtrl_logicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_shiftCtrl_valid = entries_0_uop_decoded_shiftCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_shiftCtrl_valid = io_allocateIn_payload_uop_decoded_shiftCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_shiftCtrl_isRight = entries_0_uop_decoded_shiftCtrl_isRight;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_shiftCtrl_isRight = io_allocateIn_payload_uop_decoded_shiftCtrl_isRight;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_shiftCtrl_isArithmetic = entries_0_uop_decoded_shiftCtrl_isArithmetic;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_shiftCtrl_isArithmetic = io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_shiftCtrl_isRotate = entries_0_uop_decoded_shiftCtrl_isRotate;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_shiftCtrl_isRotate = io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_shiftCtrl_isDoubleWord = entries_0_uop_decoded_shiftCtrl_isDoubleWord;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_shiftCtrl_isDoubleWord = io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_mulDivCtrl_valid = entries_0_uop_decoded_mulDivCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_mulDivCtrl_valid = io_allocateIn_payload_uop_decoded_mulDivCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_mulDivCtrl_isDiv = entries_0_uop_decoded_mulDivCtrl_isDiv;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_mulDivCtrl_isDiv = io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_mulDivCtrl_isSigned = entries_0_uop_decoded_mulDivCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_mulDivCtrl_isSigned = io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_mulDivCtrl_isWordOp = entries_0_uop_decoded_mulDivCtrl_isWordOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_mulDivCtrl_isWordOp = io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_size = entries_0_uop_decoded_memCtrl_size;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_size = io_allocateIn_payload_uop_decoded_memCtrl_size;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_isSignedLoad = entries_0_uop_decoded_memCtrl_isSignedLoad;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_isSignedLoad = io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_isStore = entries_0_uop_decoded_memCtrl_isStore;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_isStore = io_allocateIn_payload_uop_decoded_memCtrl_isStore;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_isLoadLinked = entries_0_uop_decoded_memCtrl_isLoadLinked;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_isLoadLinked = io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_isStoreCond = entries_0_uop_decoded_memCtrl_isStoreCond;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_isStoreCond = io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_atomicOp = entries_0_uop_decoded_memCtrl_atomicOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_atomicOp = io_allocateIn_payload_uop_decoded_memCtrl_atomicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_isFence = entries_0_uop_decoded_memCtrl_isFence;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_isFence = io_allocateIn_payload_uop_decoded_memCtrl_isFence;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_fenceMode = entries_0_uop_decoded_memCtrl_fenceMode;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_fenceMode = io_allocateIn_payload_uop_decoded_memCtrl_fenceMode;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_isCacheOp = entries_0_uop_decoded_memCtrl_isCacheOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_isCacheOp = io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_cacheOpType = entries_0_uop_decoded_memCtrl_cacheOpType;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_cacheOpType = io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_memCtrl_isPrefetch = entries_0_uop_decoded_memCtrl_isPrefetch;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_memCtrl_isPrefetch = io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchCtrl_condition = entries_0_uop_decoded_branchCtrl_condition;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchCtrl_condition = io_allocateIn_payload_uop_decoded_branchCtrl_condition;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchCtrl_isJump = entries_0_uop_decoded_branchCtrl_isJump;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchCtrl_isJump = io_allocateIn_payload_uop_decoded_branchCtrl_isJump;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchCtrl_isLink = entries_0_uop_decoded_branchCtrl_isLink;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchCtrl_isLink = io_allocateIn_payload_uop_decoded_branchCtrl_isLink;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchCtrl_linkReg_idx = entries_0_uop_decoded_branchCtrl_linkReg_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchCtrl_linkReg_idx = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype = entries_0_uop_decoded_branchCtrl_linkReg_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchCtrl_isIndirect = entries_0_uop_decoded_branchCtrl_isIndirect;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchCtrl_isIndirect = io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchCtrl_laCfIdx = entries_0_uop_decoded_branchCtrl_laCfIdx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchCtrl_laCfIdx = io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_opType = entries_0_uop_decoded_fpuCtrl_opType;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_opType = io_allocateIn_payload_uop_decoded_fpuCtrl_opType;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1 = entries_0_uop_decoded_fpuCtrl_fpSizeSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1 = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2 = entries_0_uop_decoded_fpuCtrl_fpSizeSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2 = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest = entries_0_uop_decoded_fpuCtrl_fpSizeDest;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_roundingMode = entries_0_uop_decoded_fpuCtrl_roundingMode;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_roundingMode = io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_isIntegerDest = entries_0_uop_decoded_fpuCtrl_isIntegerDest;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_isIntegerDest = io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_isSignedCvt = entries_0_uop_decoded_fpuCtrl_isSignedCvt;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_isSignedCvt = io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_fmaNegSrc1 = entries_0_uop_decoded_fpuCtrl_fmaNegSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_fmaNegSrc1 = io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_fpuCtrl_fcmpCond = entries_0_uop_decoded_fpuCtrl_fcmpCond;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_fpuCtrl_fcmpCond = io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_csrCtrl_csrAddr = entries_0_uop_decoded_csrCtrl_csrAddr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_csrCtrl_csrAddr = io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_csrCtrl_isWrite = entries_0_uop_decoded_csrCtrl_isWrite;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_csrCtrl_isWrite = io_allocateIn_payload_uop_decoded_csrCtrl_isWrite;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_csrCtrl_isRead = entries_0_uop_decoded_csrCtrl_isRead;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_csrCtrl_isRead = io_allocateIn_payload_uop_decoded_csrCtrl_isRead;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_csrCtrl_isExchange = entries_0_uop_decoded_csrCtrl_isExchange;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_csrCtrl_isExchange = io_allocateIn_payload_uop_decoded_csrCtrl_isExchange;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_csrCtrl_useUimmAsSrc = entries_0_uop_decoded_csrCtrl_useUimmAsSrc;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_csrCtrl_useUimmAsSrc = io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_sysCtrl_sysCode = entries_0_uop_decoded_sysCtrl_sysCode;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_sysCtrl_sysCode = io_allocateIn_payload_uop_decoded_sysCtrl_sysCode;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_sysCtrl_isExceptionReturn = entries_0_uop_decoded_sysCtrl_isExceptionReturn;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_sysCtrl_isExceptionReturn = io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_sysCtrl_isTlbOp = entries_0_uop_decoded_sysCtrl_isTlbOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_sysCtrl_isTlbOp = io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_sysCtrl_tlbOpType = entries_0_uop_decoded_sysCtrl_tlbOpType;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_sysCtrl_tlbOpType = io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_decodeExceptionCode = entries_0_uop_decoded_decodeExceptionCode;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_decodeExceptionCode = io_allocateIn_payload_uop_decoded_decodeExceptionCode;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_hasDecodeException = entries_0_uop_decoded_hasDecodeException;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_hasDecodeException = io_allocateIn_payload_uop_decoded_hasDecodeException;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_isMicrocode = entries_0_uop_decoded_isMicrocode;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_isMicrocode = io_allocateIn_payload_uop_decoded_isMicrocode;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_microcodeEntry = entries_0_uop_decoded_microcodeEntry;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_microcodeEntry = io_allocateIn_payload_uop_decoded_microcodeEntry;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_isSerializing = entries_0_uop_decoded_isSerializing;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_isSerializing = io_allocateIn_payload_uop_decoded_isSerializing;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_isBranchOrJump = entries_0_uop_decoded_isBranchOrJump;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_isBranchOrJump = io_allocateIn_payload_uop_decoded_isBranchOrJump;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchPrediction_isTaken = entries_0_uop_decoded_branchPrediction_isTaken;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchPrediction_isTaken = io_allocateIn_payload_uop_decoded_branchPrediction_isTaken;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchPrediction_target = entries_0_uop_decoded_branchPrediction_target;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchPrediction_target = io_allocateIn_payload_uop_decoded_branchPrediction_target;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_decoded_branchPrediction_wasPredicted = entries_0_uop_decoded_branchPrediction_wasPredicted;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_decoded_branchPrediction_wasPredicted = io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_physSrc1_idx = entries_0_uop_rename_physSrc1_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_physSrc1_idx = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_physSrc1IsFpr = entries_0_uop_rename_physSrc1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_physSrc1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_physSrc2_idx = entries_0_uop_rename_physSrc2_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_physSrc2_idx = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_physSrc2IsFpr = entries_0_uop_rename_physSrc2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_physSrc2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_physDest_idx = entries_0_uop_rename_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_physDestIsFpr = entries_0_uop_rename_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_oldPhysDest_idx = entries_0_uop_rename_oldPhysDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_oldPhysDest_idx = io_allocateIn_payload_uop_rename_oldPhysDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_oldPhysDestIsFpr = entries_0_uop_rename_oldPhysDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_oldPhysDestIsFpr = io_allocateIn_payload_uop_rename_oldPhysDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_allocatesPhysDest = entries_0_uop_rename_allocatesPhysDest;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_allocatesPhysDest = io_allocateIn_payload_uop_rename_allocatesPhysDest;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_rename_writesToPhysReg = entries_0_uop_rename_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_rename_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_robPtr = entries_0_uop_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_uniqueId = entries_0_uop_uniqueId;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_uniqueId = io_allocateIn_payload_uop_uniqueId;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_dispatched = entries_0_uop_dispatched;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_dispatched = io_allocateIn_payload_uop_dispatched;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_executed = entries_0_uop_executed;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_executed = io_allocateIn_payload_uop_executed;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_hasException = entries_0_uop_hasException;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_hasException = io_allocateIn_payload_uop_hasException;
      end
    end
  end

  always @(*) begin
    entriesNext_0_uop_exceptionCode = entries_0_uop_exceptionCode;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_uop_exceptionCode = io_allocateIn_payload_uop_exceptionCode;
      end
    end
  end

  always @(*) begin
    entriesNext_0_robPtr = entries_0_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_physDest_idx = entries_0_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_physDestIsFpr = entries_0_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_writesToPhysReg = entries_0_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_0_useSrc1 = entries_0_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Data = entries_0_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Tag = entries_0_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Ready = entries_0_src1Ready;
    if(when_IssueQueueComponent_l186) begin
      entriesNext_0_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_3) begin
        entriesNext_0_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1IsFpr = entries_0_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_useSrc2 = entries_0_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Data = entries_0_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Tag = entries_0_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Ready = entries_0_src2Ready;
    if(when_IssueQueueComponent_l187) begin
      entriesNext_0_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_3) begin
        entriesNext_0_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2IsFpr = entries_0_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_mulDivCtrl_valid = entries_0_mulDivCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_mulDivCtrl_valid = io_allocateIn_payload_uop_decoded_mulDivCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_0_mulDivCtrl_isDiv = entries_0_mulDivCtrl_isDiv;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_mulDivCtrl_isDiv = io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv;
      end
    end
  end

  always @(*) begin
    entriesNext_0_mulDivCtrl_isSigned = entries_0_mulDivCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_mulDivCtrl_isSigned = io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_0_mulDivCtrl_isWordOp = entries_0_mulDivCtrl_isWordOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_mulDivCtrl_isWordOp = io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_pc = entries_1_uop_decoded_pc;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_pc = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_isValid = entries_1_uop_decoded_isValid;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_isValid = io_allocateIn_payload_uop_decoded_isValid;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_uopCode = entries_1_uop_decoded_uopCode;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_uopCode = io_allocateIn_payload_uop_decoded_uopCode;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_exeUnit = entries_1_uop_decoded_exeUnit;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_exeUnit = io_allocateIn_payload_uop_decoded_exeUnit;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_isa = entries_1_uop_decoded_isa;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_isa = io_allocateIn_payload_uop_decoded_isa;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_archDest_idx = entries_1_uop_decoded_archDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_archDest_idx = io_allocateIn_payload_uop_decoded_archDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_archDest_rtype = entries_1_uop_decoded_archDest_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_archDest_rtype = io_allocateIn_payload_uop_decoded_archDest_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_writeArchDestEn = entries_1_uop_decoded_writeArchDestEn;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_writeArchDestEn = io_allocateIn_payload_uop_decoded_writeArchDestEn;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_archSrc1_idx = entries_1_uop_decoded_archSrc1_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_archSrc1_idx = io_allocateIn_payload_uop_decoded_archSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_archSrc1_rtype = entries_1_uop_decoded_archSrc1_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_archSrc1_rtype = io_allocateIn_payload_uop_decoded_archSrc1_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_useArchSrc1 = entries_1_uop_decoded_useArchSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_useArchSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_archSrc2_idx = entries_1_uop_decoded_archSrc2_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_archSrc2_idx = io_allocateIn_payload_uop_decoded_archSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_archSrc2_rtype = entries_1_uop_decoded_archSrc2_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_archSrc2_rtype = io_allocateIn_payload_uop_decoded_archSrc2_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_useArchSrc2 = entries_1_uop_decoded_useArchSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_useArchSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_usePcForAddr = entries_1_uop_decoded_usePcForAddr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_usePcForAddr = io_allocateIn_payload_uop_decoded_usePcForAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_imm = entries_1_uop_decoded_imm;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_immUsage = entries_1_uop_decoded_immUsage;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_immUsage = io_allocateIn_payload_uop_decoded_immUsage;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_aluCtrl_valid = entries_1_uop_decoded_aluCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_aluCtrl_valid = io_allocateIn_payload_uop_decoded_aluCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_aluCtrl_isSub = entries_1_uop_decoded_aluCtrl_isSub;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_aluCtrl_isSub = io_allocateIn_payload_uop_decoded_aluCtrl_isSub;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_aluCtrl_isAdd = entries_1_uop_decoded_aluCtrl_isAdd;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_aluCtrl_isAdd = io_allocateIn_payload_uop_decoded_aluCtrl_isAdd;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_aluCtrl_isSigned = entries_1_uop_decoded_aluCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_aluCtrl_isSigned = io_allocateIn_payload_uop_decoded_aluCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_aluCtrl_logicOp = entries_1_uop_decoded_aluCtrl_logicOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_aluCtrl_logicOp = io_allocateIn_payload_uop_decoded_aluCtrl_logicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_shiftCtrl_valid = entries_1_uop_decoded_shiftCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_shiftCtrl_valid = io_allocateIn_payload_uop_decoded_shiftCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_shiftCtrl_isRight = entries_1_uop_decoded_shiftCtrl_isRight;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_shiftCtrl_isRight = io_allocateIn_payload_uop_decoded_shiftCtrl_isRight;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_shiftCtrl_isArithmetic = entries_1_uop_decoded_shiftCtrl_isArithmetic;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_shiftCtrl_isArithmetic = io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_shiftCtrl_isRotate = entries_1_uop_decoded_shiftCtrl_isRotate;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_shiftCtrl_isRotate = io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_shiftCtrl_isDoubleWord = entries_1_uop_decoded_shiftCtrl_isDoubleWord;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_shiftCtrl_isDoubleWord = io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_mulDivCtrl_valid = entries_1_uop_decoded_mulDivCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_mulDivCtrl_valid = io_allocateIn_payload_uop_decoded_mulDivCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_mulDivCtrl_isDiv = entries_1_uop_decoded_mulDivCtrl_isDiv;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_mulDivCtrl_isDiv = io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_mulDivCtrl_isSigned = entries_1_uop_decoded_mulDivCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_mulDivCtrl_isSigned = io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_mulDivCtrl_isWordOp = entries_1_uop_decoded_mulDivCtrl_isWordOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_mulDivCtrl_isWordOp = io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_size = entries_1_uop_decoded_memCtrl_size;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_size = io_allocateIn_payload_uop_decoded_memCtrl_size;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_isSignedLoad = entries_1_uop_decoded_memCtrl_isSignedLoad;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_isSignedLoad = io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_isStore = entries_1_uop_decoded_memCtrl_isStore;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_isStore = io_allocateIn_payload_uop_decoded_memCtrl_isStore;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_isLoadLinked = entries_1_uop_decoded_memCtrl_isLoadLinked;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_isLoadLinked = io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_isStoreCond = entries_1_uop_decoded_memCtrl_isStoreCond;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_isStoreCond = io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_atomicOp = entries_1_uop_decoded_memCtrl_atomicOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_atomicOp = io_allocateIn_payload_uop_decoded_memCtrl_atomicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_isFence = entries_1_uop_decoded_memCtrl_isFence;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_isFence = io_allocateIn_payload_uop_decoded_memCtrl_isFence;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_fenceMode = entries_1_uop_decoded_memCtrl_fenceMode;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_fenceMode = io_allocateIn_payload_uop_decoded_memCtrl_fenceMode;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_isCacheOp = entries_1_uop_decoded_memCtrl_isCacheOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_isCacheOp = io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_cacheOpType = entries_1_uop_decoded_memCtrl_cacheOpType;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_cacheOpType = io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_memCtrl_isPrefetch = entries_1_uop_decoded_memCtrl_isPrefetch;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_memCtrl_isPrefetch = io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchCtrl_condition = entries_1_uop_decoded_branchCtrl_condition;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchCtrl_condition = io_allocateIn_payload_uop_decoded_branchCtrl_condition;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchCtrl_isJump = entries_1_uop_decoded_branchCtrl_isJump;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchCtrl_isJump = io_allocateIn_payload_uop_decoded_branchCtrl_isJump;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchCtrl_isLink = entries_1_uop_decoded_branchCtrl_isLink;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchCtrl_isLink = io_allocateIn_payload_uop_decoded_branchCtrl_isLink;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchCtrl_linkReg_idx = entries_1_uop_decoded_branchCtrl_linkReg_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchCtrl_linkReg_idx = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype = entries_1_uop_decoded_branchCtrl_linkReg_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchCtrl_isIndirect = entries_1_uop_decoded_branchCtrl_isIndirect;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchCtrl_isIndirect = io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchCtrl_laCfIdx = entries_1_uop_decoded_branchCtrl_laCfIdx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchCtrl_laCfIdx = io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_opType = entries_1_uop_decoded_fpuCtrl_opType;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_opType = io_allocateIn_payload_uop_decoded_fpuCtrl_opType;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1 = entries_1_uop_decoded_fpuCtrl_fpSizeSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1 = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2 = entries_1_uop_decoded_fpuCtrl_fpSizeSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2 = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest = entries_1_uop_decoded_fpuCtrl_fpSizeDest;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_roundingMode = entries_1_uop_decoded_fpuCtrl_roundingMode;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_roundingMode = io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_isIntegerDest = entries_1_uop_decoded_fpuCtrl_isIntegerDest;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_isIntegerDest = io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_isSignedCvt = entries_1_uop_decoded_fpuCtrl_isSignedCvt;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_isSignedCvt = io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_fmaNegSrc1 = entries_1_uop_decoded_fpuCtrl_fmaNegSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_fmaNegSrc1 = io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_fpuCtrl_fcmpCond = entries_1_uop_decoded_fpuCtrl_fcmpCond;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_fpuCtrl_fcmpCond = io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_csrCtrl_csrAddr = entries_1_uop_decoded_csrCtrl_csrAddr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_csrCtrl_csrAddr = io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_csrCtrl_isWrite = entries_1_uop_decoded_csrCtrl_isWrite;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_csrCtrl_isWrite = io_allocateIn_payload_uop_decoded_csrCtrl_isWrite;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_csrCtrl_isRead = entries_1_uop_decoded_csrCtrl_isRead;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_csrCtrl_isRead = io_allocateIn_payload_uop_decoded_csrCtrl_isRead;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_csrCtrl_isExchange = entries_1_uop_decoded_csrCtrl_isExchange;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_csrCtrl_isExchange = io_allocateIn_payload_uop_decoded_csrCtrl_isExchange;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_csrCtrl_useUimmAsSrc = entries_1_uop_decoded_csrCtrl_useUimmAsSrc;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_csrCtrl_useUimmAsSrc = io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_sysCtrl_sysCode = entries_1_uop_decoded_sysCtrl_sysCode;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_sysCtrl_sysCode = io_allocateIn_payload_uop_decoded_sysCtrl_sysCode;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_sysCtrl_isExceptionReturn = entries_1_uop_decoded_sysCtrl_isExceptionReturn;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_sysCtrl_isExceptionReturn = io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_sysCtrl_isTlbOp = entries_1_uop_decoded_sysCtrl_isTlbOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_sysCtrl_isTlbOp = io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_sysCtrl_tlbOpType = entries_1_uop_decoded_sysCtrl_tlbOpType;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_sysCtrl_tlbOpType = io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_decodeExceptionCode = entries_1_uop_decoded_decodeExceptionCode;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_decodeExceptionCode = io_allocateIn_payload_uop_decoded_decodeExceptionCode;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_hasDecodeException = entries_1_uop_decoded_hasDecodeException;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_hasDecodeException = io_allocateIn_payload_uop_decoded_hasDecodeException;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_isMicrocode = entries_1_uop_decoded_isMicrocode;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_isMicrocode = io_allocateIn_payload_uop_decoded_isMicrocode;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_microcodeEntry = entries_1_uop_decoded_microcodeEntry;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_microcodeEntry = io_allocateIn_payload_uop_decoded_microcodeEntry;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_isSerializing = entries_1_uop_decoded_isSerializing;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_isSerializing = io_allocateIn_payload_uop_decoded_isSerializing;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_isBranchOrJump = entries_1_uop_decoded_isBranchOrJump;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_isBranchOrJump = io_allocateIn_payload_uop_decoded_isBranchOrJump;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchPrediction_isTaken = entries_1_uop_decoded_branchPrediction_isTaken;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchPrediction_isTaken = io_allocateIn_payload_uop_decoded_branchPrediction_isTaken;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchPrediction_target = entries_1_uop_decoded_branchPrediction_target;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchPrediction_target = io_allocateIn_payload_uop_decoded_branchPrediction_target;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_decoded_branchPrediction_wasPredicted = entries_1_uop_decoded_branchPrediction_wasPredicted;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_decoded_branchPrediction_wasPredicted = io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_physSrc1_idx = entries_1_uop_rename_physSrc1_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_physSrc1_idx = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_physSrc1IsFpr = entries_1_uop_rename_physSrc1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_physSrc1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_physSrc2_idx = entries_1_uop_rename_physSrc2_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_physSrc2_idx = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_physSrc2IsFpr = entries_1_uop_rename_physSrc2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_physSrc2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_physDest_idx = entries_1_uop_rename_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_physDestIsFpr = entries_1_uop_rename_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_oldPhysDest_idx = entries_1_uop_rename_oldPhysDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_oldPhysDest_idx = io_allocateIn_payload_uop_rename_oldPhysDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_oldPhysDestIsFpr = entries_1_uop_rename_oldPhysDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_oldPhysDestIsFpr = io_allocateIn_payload_uop_rename_oldPhysDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_allocatesPhysDest = entries_1_uop_rename_allocatesPhysDest;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_allocatesPhysDest = io_allocateIn_payload_uop_rename_allocatesPhysDest;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_rename_writesToPhysReg = entries_1_uop_rename_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_rename_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_robPtr = entries_1_uop_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_uniqueId = entries_1_uop_uniqueId;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_uniqueId = io_allocateIn_payload_uop_uniqueId;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_dispatched = entries_1_uop_dispatched;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_dispatched = io_allocateIn_payload_uop_dispatched;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_executed = entries_1_uop_executed;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_executed = io_allocateIn_payload_uop_executed;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_hasException = entries_1_uop_hasException;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_hasException = io_allocateIn_payload_uop_hasException;
      end
    end
  end

  always @(*) begin
    entriesNext_1_uop_exceptionCode = entries_1_uop_exceptionCode;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_uop_exceptionCode = io_allocateIn_payload_uop_exceptionCode;
      end
    end
  end

  always @(*) begin
    entriesNext_1_robPtr = entries_1_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_physDest_idx = entries_1_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_physDestIsFpr = entries_1_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_writesToPhysReg = entries_1_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_1_useSrc1 = entries_1_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Data = entries_1_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Tag = entries_1_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Ready = entries_1_src1Ready;
    if(when_IssueQueueComponent_l186_1) begin
      entriesNext_1_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_4) begin
        entriesNext_1_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1IsFpr = entries_1_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_useSrc2 = entries_1_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Data = entries_1_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Tag = entries_1_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Ready = entries_1_src2Ready;
    if(when_IssueQueueComponent_l187_1) begin
      entriesNext_1_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_4) begin
        entriesNext_1_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2IsFpr = entries_1_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_mulDivCtrl_valid = entries_1_mulDivCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_mulDivCtrl_valid = io_allocateIn_payload_uop_decoded_mulDivCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_1_mulDivCtrl_isDiv = entries_1_mulDivCtrl_isDiv;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_mulDivCtrl_isDiv = io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv;
      end
    end
  end

  always @(*) begin
    entriesNext_1_mulDivCtrl_isSigned = entries_1_mulDivCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_mulDivCtrl_isSigned = io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_1_mulDivCtrl_isWordOp = entries_1_mulDivCtrl_isWordOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_mulDivCtrl_isWordOp = io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_pc = entries_2_uop_decoded_pc;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_pc = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_isValid = entries_2_uop_decoded_isValid;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_isValid = io_allocateIn_payload_uop_decoded_isValid;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_uopCode = entries_2_uop_decoded_uopCode;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_uopCode = io_allocateIn_payload_uop_decoded_uopCode;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_exeUnit = entries_2_uop_decoded_exeUnit;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_exeUnit = io_allocateIn_payload_uop_decoded_exeUnit;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_isa = entries_2_uop_decoded_isa;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_isa = io_allocateIn_payload_uop_decoded_isa;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_archDest_idx = entries_2_uop_decoded_archDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_archDest_idx = io_allocateIn_payload_uop_decoded_archDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_archDest_rtype = entries_2_uop_decoded_archDest_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_archDest_rtype = io_allocateIn_payload_uop_decoded_archDest_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_writeArchDestEn = entries_2_uop_decoded_writeArchDestEn;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_writeArchDestEn = io_allocateIn_payload_uop_decoded_writeArchDestEn;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_archSrc1_idx = entries_2_uop_decoded_archSrc1_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_archSrc1_idx = io_allocateIn_payload_uop_decoded_archSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_archSrc1_rtype = entries_2_uop_decoded_archSrc1_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_archSrc1_rtype = io_allocateIn_payload_uop_decoded_archSrc1_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_useArchSrc1 = entries_2_uop_decoded_useArchSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_useArchSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_archSrc2_idx = entries_2_uop_decoded_archSrc2_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_archSrc2_idx = io_allocateIn_payload_uop_decoded_archSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_archSrc2_rtype = entries_2_uop_decoded_archSrc2_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_archSrc2_rtype = io_allocateIn_payload_uop_decoded_archSrc2_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_useArchSrc2 = entries_2_uop_decoded_useArchSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_useArchSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_usePcForAddr = entries_2_uop_decoded_usePcForAddr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_usePcForAddr = io_allocateIn_payload_uop_decoded_usePcForAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_imm = entries_2_uop_decoded_imm;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_immUsage = entries_2_uop_decoded_immUsage;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_immUsage = io_allocateIn_payload_uop_decoded_immUsage;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_aluCtrl_valid = entries_2_uop_decoded_aluCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_aluCtrl_valid = io_allocateIn_payload_uop_decoded_aluCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_aluCtrl_isSub = entries_2_uop_decoded_aluCtrl_isSub;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_aluCtrl_isSub = io_allocateIn_payload_uop_decoded_aluCtrl_isSub;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_aluCtrl_isAdd = entries_2_uop_decoded_aluCtrl_isAdd;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_aluCtrl_isAdd = io_allocateIn_payload_uop_decoded_aluCtrl_isAdd;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_aluCtrl_isSigned = entries_2_uop_decoded_aluCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_aluCtrl_isSigned = io_allocateIn_payload_uop_decoded_aluCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_aluCtrl_logicOp = entries_2_uop_decoded_aluCtrl_logicOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_aluCtrl_logicOp = io_allocateIn_payload_uop_decoded_aluCtrl_logicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_shiftCtrl_valid = entries_2_uop_decoded_shiftCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_shiftCtrl_valid = io_allocateIn_payload_uop_decoded_shiftCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_shiftCtrl_isRight = entries_2_uop_decoded_shiftCtrl_isRight;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_shiftCtrl_isRight = io_allocateIn_payload_uop_decoded_shiftCtrl_isRight;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_shiftCtrl_isArithmetic = entries_2_uop_decoded_shiftCtrl_isArithmetic;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_shiftCtrl_isArithmetic = io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_shiftCtrl_isRotate = entries_2_uop_decoded_shiftCtrl_isRotate;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_shiftCtrl_isRotate = io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_shiftCtrl_isDoubleWord = entries_2_uop_decoded_shiftCtrl_isDoubleWord;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_shiftCtrl_isDoubleWord = io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_mulDivCtrl_valid = entries_2_uop_decoded_mulDivCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_mulDivCtrl_valid = io_allocateIn_payload_uop_decoded_mulDivCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_mulDivCtrl_isDiv = entries_2_uop_decoded_mulDivCtrl_isDiv;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_mulDivCtrl_isDiv = io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_mulDivCtrl_isSigned = entries_2_uop_decoded_mulDivCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_mulDivCtrl_isSigned = io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_mulDivCtrl_isWordOp = entries_2_uop_decoded_mulDivCtrl_isWordOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_mulDivCtrl_isWordOp = io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_size = entries_2_uop_decoded_memCtrl_size;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_size = io_allocateIn_payload_uop_decoded_memCtrl_size;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_isSignedLoad = entries_2_uop_decoded_memCtrl_isSignedLoad;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_isSignedLoad = io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_isStore = entries_2_uop_decoded_memCtrl_isStore;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_isStore = io_allocateIn_payload_uop_decoded_memCtrl_isStore;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_isLoadLinked = entries_2_uop_decoded_memCtrl_isLoadLinked;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_isLoadLinked = io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_isStoreCond = entries_2_uop_decoded_memCtrl_isStoreCond;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_isStoreCond = io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_atomicOp = entries_2_uop_decoded_memCtrl_atomicOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_atomicOp = io_allocateIn_payload_uop_decoded_memCtrl_atomicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_isFence = entries_2_uop_decoded_memCtrl_isFence;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_isFence = io_allocateIn_payload_uop_decoded_memCtrl_isFence;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_fenceMode = entries_2_uop_decoded_memCtrl_fenceMode;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_fenceMode = io_allocateIn_payload_uop_decoded_memCtrl_fenceMode;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_isCacheOp = entries_2_uop_decoded_memCtrl_isCacheOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_isCacheOp = io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_cacheOpType = entries_2_uop_decoded_memCtrl_cacheOpType;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_cacheOpType = io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_memCtrl_isPrefetch = entries_2_uop_decoded_memCtrl_isPrefetch;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_memCtrl_isPrefetch = io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchCtrl_condition = entries_2_uop_decoded_branchCtrl_condition;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchCtrl_condition = io_allocateIn_payload_uop_decoded_branchCtrl_condition;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchCtrl_isJump = entries_2_uop_decoded_branchCtrl_isJump;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchCtrl_isJump = io_allocateIn_payload_uop_decoded_branchCtrl_isJump;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchCtrl_isLink = entries_2_uop_decoded_branchCtrl_isLink;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchCtrl_isLink = io_allocateIn_payload_uop_decoded_branchCtrl_isLink;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchCtrl_linkReg_idx = entries_2_uop_decoded_branchCtrl_linkReg_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchCtrl_linkReg_idx = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype = entries_2_uop_decoded_branchCtrl_linkReg_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchCtrl_isIndirect = entries_2_uop_decoded_branchCtrl_isIndirect;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchCtrl_isIndirect = io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchCtrl_laCfIdx = entries_2_uop_decoded_branchCtrl_laCfIdx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchCtrl_laCfIdx = io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_opType = entries_2_uop_decoded_fpuCtrl_opType;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_opType = io_allocateIn_payload_uop_decoded_fpuCtrl_opType;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1 = entries_2_uop_decoded_fpuCtrl_fpSizeSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1 = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2 = entries_2_uop_decoded_fpuCtrl_fpSizeSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2 = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest = entries_2_uop_decoded_fpuCtrl_fpSizeDest;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_roundingMode = entries_2_uop_decoded_fpuCtrl_roundingMode;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_roundingMode = io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_isIntegerDest = entries_2_uop_decoded_fpuCtrl_isIntegerDest;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_isIntegerDest = io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_isSignedCvt = entries_2_uop_decoded_fpuCtrl_isSignedCvt;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_isSignedCvt = io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_fmaNegSrc1 = entries_2_uop_decoded_fpuCtrl_fmaNegSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_fmaNegSrc1 = io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_fpuCtrl_fcmpCond = entries_2_uop_decoded_fpuCtrl_fcmpCond;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_fpuCtrl_fcmpCond = io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_csrCtrl_csrAddr = entries_2_uop_decoded_csrCtrl_csrAddr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_csrCtrl_csrAddr = io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_csrCtrl_isWrite = entries_2_uop_decoded_csrCtrl_isWrite;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_csrCtrl_isWrite = io_allocateIn_payload_uop_decoded_csrCtrl_isWrite;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_csrCtrl_isRead = entries_2_uop_decoded_csrCtrl_isRead;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_csrCtrl_isRead = io_allocateIn_payload_uop_decoded_csrCtrl_isRead;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_csrCtrl_isExchange = entries_2_uop_decoded_csrCtrl_isExchange;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_csrCtrl_isExchange = io_allocateIn_payload_uop_decoded_csrCtrl_isExchange;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_csrCtrl_useUimmAsSrc = entries_2_uop_decoded_csrCtrl_useUimmAsSrc;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_csrCtrl_useUimmAsSrc = io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_sysCtrl_sysCode = entries_2_uop_decoded_sysCtrl_sysCode;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_sysCtrl_sysCode = io_allocateIn_payload_uop_decoded_sysCtrl_sysCode;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_sysCtrl_isExceptionReturn = entries_2_uop_decoded_sysCtrl_isExceptionReturn;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_sysCtrl_isExceptionReturn = io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_sysCtrl_isTlbOp = entries_2_uop_decoded_sysCtrl_isTlbOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_sysCtrl_isTlbOp = io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_sysCtrl_tlbOpType = entries_2_uop_decoded_sysCtrl_tlbOpType;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_sysCtrl_tlbOpType = io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_decodeExceptionCode = entries_2_uop_decoded_decodeExceptionCode;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_decodeExceptionCode = io_allocateIn_payload_uop_decoded_decodeExceptionCode;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_hasDecodeException = entries_2_uop_decoded_hasDecodeException;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_hasDecodeException = io_allocateIn_payload_uop_decoded_hasDecodeException;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_isMicrocode = entries_2_uop_decoded_isMicrocode;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_isMicrocode = io_allocateIn_payload_uop_decoded_isMicrocode;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_microcodeEntry = entries_2_uop_decoded_microcodeEntry;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_microcodeEntry = io_allocateIn_payload_uop_decoded_microcodeEntry;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_isSerializing = entries_2_uop_decoded_isSerializing;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_isSerializing = io_allocateIn_payload_uop_decoded_isSerializing;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_isBranchOrJump = entries_2_uop_decoded_isBranchOrJump;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_isBranchOrJump = io_allocateIn_payload_uop_decoded_isBranchOrJump;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchPrediction_isTaken = entries_2_uop_decoded_branchPrediction_isTaken;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchPrediction_isTaken = io_allocateIn_payload_uop_decoded_branchPrediction_isTaken;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchPrediction_target = entries_2_uop_decoded_branchPrediction_target;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchPrediction_target = io_allocateIn_payload_uop_decoded_branchPrediction_target;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_decoded_branchPrediction_wasPredicted = entries_2_uop_decoded_branchPrediction_wasPredicted;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_decoded_branchPrediction_wasPredicted = io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_physSrc1_idx = entries_2_uop_rename_physSrc1_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_physSrc1_idx = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_physSrc1IsFpr = entries_2_uop_rename_physSrc1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_physSrc1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_physSrc2_idx = entries_2_uop_rename_physSrc2_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_physSrc2_idx = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_physSrc2IsFpr = entries_2_uop_rename_physSrc2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_physSrc2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_physDest_idx = entries_2_uop_rename_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_physDestIsFpr = entries_2_uop_rename_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_oldPhysDest_idx = entries_2_uop_rename_oldPhysDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_oldPhysDest_idx = io_allocateIn_payload_uop_rename_oldPhysDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_oldPhysDestIsFpr = entries_2_uop_rename_oldPhysDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_oldPhysDestIsFpr = io_allocateIn_payload_uop_rename_oldPhysDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_allocatesPhysDest = entries_2_uop_rename_allocatesPhysDest;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_allocatesPhysDest = io_allocateIn_payload_uop_rename_allocatesPhysDest;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_rename_writesToPhysReg = entries_2_uop_rename_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_rename_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_robPtr = entries_2_uop_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_uniqueId = entries_2_uop_uniqueId;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_uniqueId = io_allocateIn_payload_uop_uniqueId;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_dispatched = entries_2_uop_dispatched;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_dispatched = io_allocateIn_payload_uop_dispatched;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_executed = entries_2_uop_executed;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_executed = io_allocateIn_payload_uop_executed;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_hasException = entries_2_uop_hasException;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_hasException = io_allocateIn_payload_uop_hasException;
      end
    end
  end

  always @(*) begin
    entriesNext_2_uop_exceptionCode = entries_2_uop_exceptionCode;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_uop_exceptionCode = io_allocateIn_payload_uop_exceptionCode;
      end
    end
  end

  always @(*) begin
    entriesNext_2_robPtr = entries_2_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_physDest_idx = entries_2_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_physDestIsFpr = entries_2_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_writesToPhysReg = entries_2_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_2_useSrc1 = entries_2_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Data = entries_2_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Tag = entries_2_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Ready = entries_2_src1Ready;
    if(when_IssueQueueComponent_l186_2) begin
      entriesNext_2_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_5) begin
        entriesNext_2_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1IsFpr = entries_2_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_useSrc2 = entries_2_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Data = entries_2_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Tag = entries_2_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Ready = entries_2_src2Ready;
    if(when_IssueQueueComponent_l187_2) begin
      entriesNext_2_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_5) begin
        entriesNext_2_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2IsFpr = entries_2_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_mulDivCtrl_valid = entries_2_mulDivCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_mulDivCtrl_valid = io_allocateIn_payload_uop_decoded_mulDivCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_2_mulDivCtrl_isDiv = entries_2_mulDivCtrl_isDiv;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_mulDivCtrl_isDiv = io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv;
      end
    end
  end

  always @(*) begin
    entriesNext_2_mulDivCtrl_isSigned = entries_2_mulDivCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_mulDivCtrl_isSigned = io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_2_mulDivCtrl_isWordOp = entries_2_mulDivCtrl_isWordOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_mulDivCtrl_isWordOp = io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_pc = entries_3_uop_decoded_pc;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_pc = io_allocateIn_payload_uop_decoded_pc;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_isValid = entries_3_uop_decoded_isValid;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_isValid = io_allocateIn_payload_uop_decoded_isValid;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_uopCode = entries_3_uop_decoded_uopCode;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_uopCode = io_allocateIn_payload_uop_decoded_uopCode;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_exeUnit = entries_3_uop_decoded_exeUnit;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_exeUnit = io_allocateIn_payload_uop_decoded_exeUnit;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_isa = entries_3_uop_decoded_isa;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_isa = io_allocateIn_payload_uop_decoded_isa;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_archDest_idx = entries_3_uop_decoded_archDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_archDest_idx = io_allocateIn_payload_uop_decoded_archDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_archDest_rtype = entries_3_uop_decoded_archDest_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_archDest_rtype = io_allocateIn_payload_uop_decoded_archDest_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_writeArchDestEn = entries_3_uop_decoded_writeArchDestEn;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_writeArchDestEn = io_allocateIn_payload_uop_decoded_writeArchDestEn;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_archSrc1_idx = entries_3_uop_decoded_archSrc1_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_archSrc1_idx = io_allocateIn_payload_uop_decoded_archSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_archSrc1_rtype = entries_3_uop_decoded_archSrc1_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_archSrc1_rtype = io_allocateIn_payload_uop_decoded_archSrc1_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_useArchSrc1 = entries_3_uop_decoded_useArchSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_useArchSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_archSrc2_idx = entries_3_uop_decoded_archSrc2_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_archSrc2_idx = io_allocateIn_payload_uop_decoded_archSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_archSrc2_rtype = entries_3_uop_decoded_archSrc2_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_archSrc2_rtype = io_allocateIn_payload_uop_decoded_archSrc2_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_useArchSrc2 = entries_3_uop_decoded_useArchSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_useArchSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_usePcForAddr = entries_3_uop_decoded_usePcForAddr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_usePcForAddr = io_allocateIn_payload_uop_decoded_usePcForAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_imm = entries_3_uop_decoded_imm;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_immUsage = entries_3_uop_decoded_immUsage;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_immUsage = io_allocateIn_payload_uop_decoded_immUsage;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_aluCtrl_valid = entries_3_uop_decoded_aluCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_aluCtrl_valid = io_allocateIn_payload_uop_decoded_aluCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_aluCtrl_isSub = entries_3_uop_decoded_aluCtrl_isSub;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_aluCtrl_isSub = io_allocateIn_payload_uop_decoded_aluCtrl_isSub;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_aluCtrl_isAdd = entries_3_uop_decoded_aluCtrl_isAdd;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_aluCtrl_isAdd = io_allocateIn_payload_uop_decoded_aluCtrl_isAdd;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_aluCtrl_isSigned = entries_3_uop_decoded_aluCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_aluCtrl_isSigned = io_allocateIn_payload_uop_decoded_aluCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_aluCtrl_logicOp = entries_3_uop_decoded_aluCtrl_logicOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_aluCtrl_logicOp = io_allocateIn_payload_uop_decoded_aluCtrl_logicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_shiftCtrl_valid = entries_3_uop_decoded_shiftCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_shiftCtrl_valid = io_allocateIn_payload_uop_decoded_shiftCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_shiftCtrl_isRight = entries_3_uop_decoded_shiftCtrl_isRight;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_shiftCtrl_isRight = io_allocateIn_payload_uop_decoded_shiftCtrl_isRight;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_shiftCtrl_isArithmetic = entries_3_uop_decoded_shiftCtrl_isArithmetic;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_shiftCtrl_isArithmetic = io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_shiftCtrl_isRotate = entries_3_uop_decoded_shiftCtrl_isRotate;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_shiftCtrl_isRotate = io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_shiftCtrl_isDoubleWord = entries_3_uop_decoded_shiftCtrl_isDoubleWord;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_shiftCtrl_isDoubleWord = io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_mulDivCtrl_valid = entries_3_uop_decoded_mulDivCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_mulDivCtrl_valid = io_allocateIn_payload_uop_decoded_mulDivCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_mulDivCtrl_isDiv = entries_3_uop_decoded_mulDivCtrl_isDiv;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_mulDivCtrl_isDiv = io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_mulDivCtrl_isSigned = entries_3_uop_decoded_mulDivCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_mulDivCtrl_isSigned = io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_mulDivCtrl_isWordOp = entries_3_uop_decoded_mulDivCtrl_isWordOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_mulDivCtrl_isWordOp = io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_size = entries_3_uop_decoded_memCtrl_size;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_size = io_allocateIn_payload_uop_decoded_memCtrl_size;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_isSignedLoad = entries_3_uop_decoded_memCtrl_isSignedLoad;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_isSignedLoad = io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_isStore = entries_3_uop_decoded_memCtrl_isStore;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_isStore = io_allocateIn_payload_uop_decoded_memCtrl_isStore;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_isLoadLinked = entries_3_uop_decoded_memCtrl_isLoadLinked;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_isLoadLinked = io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_isStoreCond = entries_3_uop_decoded_memCtrl_isStoreCond;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_isStoreCond = io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_atomicOp = entries_3_uop_decoded_memCtrl_atomicOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_atomicOp = io_allocateIn_payload_uop_decoded_memCtrl_atomicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_isFence = entries_3_uop_decoded_memCtrl_isFence;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_isFence = io_allocateIn_payload_uop_decoded_memCtrl_isFence;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_fenceMode = entries_3_uop_decoded_memCtrl_fenceMode;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_fenceMode = io_allocateIn_payload_uop_decoded_memCtrl_fenceMode;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_isCacheOp = entries_3_uop_decoded_memCtrl_isCacheOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_isCacheOp = io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_cacheOpType = entries_3_uop_decoded_memCtrl_cacheOpType;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_cacheOpType = io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_memCtrl_isPrefetch = entries_3_uop_decoded_memCtrl_isPrefetch;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_memCtrl_isPrefetch = io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchCtrl_condition = entries_3_uop_decoded_branchCtrl_condition;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchCtrl_condition = io_allocateIn_payload_uop_decoded_branchCtrl_condition;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchCtrl_isJump = entries_3_uop_decoded_branchCtrl_isJump;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchCtrl_isJump = io_allocateIn_payload_uop_decoded_branchCtrl_isJump;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchCtrl_isLink = entries_3_uop_decoded_branchCtrl_isLink;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchCtrl_isLink = io_allocateIn_payload_uop_decoded_branchCtrl_isLink;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchCtrl_linkReg_idx = entries_3_uop_decoded_branchCtrl_linkReg_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchCtrl_linkReg_idx = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype = entries_3_uop_decoded_branchCtrl_linkReg_rtype;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype = io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchCtrl_isIndirect = entries_3_uop_decoded_branchCtrl_isIndirect;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchCtrl_isIndirect = io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchCtrl_laCfIdx = entries_3_uop_decoded_branchCtrl_laCfIdx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchCtrl_laCfIdx = io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_opType = entries_3_uop_decoded_fpuCtrl_opType;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_opType = io_allocateIn_payload_uop_decoded_fpuCtrl_opType;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1 = entries_3_uop_decoded_fpuCtrl_fpSizeSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1 = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2 = entries_3_uop_decoded_fpuCtrl_fpSizeSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2 = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest = entries_3_uop_decoded_fpuCtrl_fpSizeDest;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest = io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_roundingMode = entries_3_uop_decoded_fpuCtrl_roundingMode;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_roundingMode = io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_isIntegerDest = entries_3_uop_decoded_fpuCtrl_isIntegerDest;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_isIntegerDest = io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_isSignedCvt = entries_3_uop_decoded_fpuCtrl_isSignedCvt;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_isSignedCvt = io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_fmaNegSrc1 = entries_3_uop_decoded_fpuCtrl_fmaNegSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_fmaNegSrc1 = io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_fpuCtrl_fcmpCond = entries_3_uop_decoded_fpuCtrl_fcmpCond;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_fpuCtrl_fcmpCond = io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_csrCtrl_csrAddr = entries_3_uop_decoded_csrCtrl_csrAddr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_csrCtrl_csrAddr = io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_csrCtrl_isWrite = entries_3_uop_decoded_csrCtrl_isWrite;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_csrCtrl_isWrite = io_allocateIn_payload_uop_decoded_csrCtrl_isWrite;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_csrCtrl_isRead = entries_3_uop_decoded_csrCtrl_isRead;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_csrCtrl_isRead = io_allocateIn_payload_uop_decoded_csrCtrl_isRead;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_csrCtrl_isExchange = entries_3_uop_decoded_csrCtrl_isExchange;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_csrCtrl_isExchange = io_allocateIn_payload_uop_decoded_csrCtrl_isExchange;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_csrCtrl_useUimmAsSrc = entries_3_uop_decoded_csrCtrl_useUimmAsSrc;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_csrCtrl_useUimmAsSrc = io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_sysCtrl_sysCode = entries_3_uop_decoded_sysCtrl_sysCode;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_sysCtrl_sysCode = io_allocateIn_payload_uop_decoded_sysCtrl_sysCode;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_sysCtrl_isExceptionReturn = entries_3_uop_decoded_sysCtrl_isExceptionReturn;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_sysCtrl_isExceptionReturn = io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_sysCtrl_isTlbOp = entries_3_uop_decoded_sysCtrl_isTlbOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_sysCtrl_isTlbOp = io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_sysCtrl_tlbOpType = entries_3_uop_decoded_sysCtrl_tlbOpType;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_sysCtrl_tlbOpType = io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_decodeExceptionCode = entries_3_uop_decoded_decodeExceptionCode;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_decodeExceptionCode = io_allocateIn_payload_uop_decoded_decodeExceptionCode;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_hasDecodeException = entries_3_uop_decoded_hasDecodeException;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_hasDecodeException = io_allocateIn_payload_uop_decoded_hasDecodeException;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_isMicrocode = entries_3_uop_decoded_isMicrocode;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_isMicrocode = io_allocateIn_payload_uop_decoded_isMicrocode;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_microcodeEntry = entries_3_uop_decoded_microcodeEntry;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_microcodeEntry = io_allocateIn_payload_uop_decoded_microcodeEntry;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_isSerializing = entries_3_uop_decoded_isSerializing;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_isSerializing = io_allocateIn_payload_uop_decoded_isSerializing;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_isBranchOrJump = entries_3_uop_decoded_isBranchOrJump;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_isBranchOrJump = io_allocateIn_payload_uop_decoded_isBranchOrJump;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchPrediction_isTaken = entries_3_uop_decoded_branchPrediction_isTaken;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchPrediction_isTaken = io_allocateIn_payload_uop_decoded_branchPrediction_isTaken;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchPrediction_target = entries_3_uop_decoded_branchPrediction_target;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchPrediction_target = io_allocateIn_payload_uop_decoded_branchPrediction_target;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_decoded_branchPrediction_wasPredicted = entries_3_uop_decoded_branchPrediction_wasPredicted;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_decoded_branchPrediction_wasPredicted = io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_physSrc1_idx = entries_3_uop_rename_physSrc1_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_physSrc1_idx = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_physSrc1IsFpr = entries_3_uop_rename_physSrc1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_physSrc1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_physSrc2_idx = entries_3_uop_rename_physSrc2_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_physSrc2_idx = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_physSrc2IsFpr = entries_3_uop_rename_physSrc2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_physSrc2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_physDest_idx = entries_3_uop_rename_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_physDestIsFpr = entries_3_uop_rename_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_oldPhysDest_idx = entries_3_uop_rename_oldPhysDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_oldPhysDest_idx = io_allocateIn_payload_uop_rename_oldPhysDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_oldPhysDestIsFpr = entries_3_uop_rename_oldPhysDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_oldPhysDestIsFpr = io_allocateIn_payload_uop_rename_oldPhysDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_allocatesPhysDest = entries_3_uop_rename_allocatesPhysDest;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_allocatesPhysDest = io_allocateIn_payload_uop_rename_allocatesPhysDest;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_rename_writesToPhysReg = entries_3_uop_rename_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_rename_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_robPtr = entries_3_uop_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_uniqueId = entries_3_uop_uniqueId;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_uniqueId = io_allocateIn_payload_uop_uniqueId;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_dispatched = entries_3_uop_dispatched;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_dispatched = io_allocateIn_payload_uop_dispatched;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_executed = entries_3_uop_executed;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_executed = io_allocateIn_payload_uop_executed;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_hasException = entries_3_uop_hasException;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_hasException = io_allocateIn_payload_uop_hasException;
      end
    end
  end

  always @(*) begin
    entriesNext_3_uop_exceptionCode = entries_3_uop_exceptionCode;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_uop_exceptionCode = io_allocateIn_payload_uop_exceptionCode;
      end
    end
  end

  always @(*) begin
    entriesNext_3_robPtr = entries_3_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_physDest_idx = entries_3_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_physDestIsFpr = entries_3_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_writesToPhysReg = entries_3_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_3_useSrc1 = entries_3_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Data = entries_3_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Tag = entries_3_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Ready = entries_3_src1Ready;
    if(when_IssueQueueComponent_l186_3) begin
      entriesNext_3_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_6) begin
        entriesNext_3_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1IsFpr = entries_3_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_useSrc2 = entries_3_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Data = entries_3_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Tag = entries_3_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Ready = entries_3_src2Ready;
    if(when_IssueQueueComponent_l187_3) begin
      entriesNext_3_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_6) begin
        entriesNext_3_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2IsFpr = entries_3_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_mulDivCtrl_valid = entries_3_mulDivCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_mulDivCtrl_valid = io_allocateIn_payload_uop_decoded_mulDivCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_3_mulDivCtrl_isDiv = entries_3_mulDivCtrl_isDiv;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_mulDivCtrl_isDiv = io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv;
      end
    end
  end

  always @(*) begin
    entriesNext_3_mulDivCtrl_isSigned = entries_3_mulDivCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_mulDivCtrl_isSigned = io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_3_mulDivCtrl_isWordOp = entries_3_mulDivCtrl_isWordOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_mulDivCtrl_isWordOp = io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp;
      end
    end
  end

  always @(*) begin
    entryValidsNext_0 = entryValids_0;
    if(io_issueOut_fire) begin
      if(_zz_1[0]) begin
        entryValidsNext_0 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[0]) begin
        entryValidsNext_0 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_0 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_1 = entryValids_1;
    if(io_issueOut_fire) begin
      if(_zz_1[1]) begin
        entryValidsNext_1 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[1]) begin
        entryValidsNext_1 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_1 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_2 = entryValids_2;
    if(io_issueOut_fire) begin
      if(_zz_1[2]) begin
        entryValidsNext_2 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[2]) begin
        entryValidsNext_2 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_2 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_3 = entryValids_3;
    if(io_issueOut_fire) begin
      if(_zz_1[3]) begin
        entryValidsNext_3 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[3]) begin
        entryValidsNext_3 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_3 = 1'b0;
    end
  end

  assign when_IssueQueueComponent_l186 = wokeUpSrc1Mask[0];
  assign when_IssueQueueComponent_l187 = wokeUpSrc2Mask[0];
  assign when_IssueQueueComponent_l186_1 = wokeUpSrc1Mask[1];
  assign when_IssueQueueComponent_l187_1 = wokeUpSrc2Mask[1];
  assign when_IssueQueueComponent_l186_2 = wokeUpSrc1Mask[2];
  assign when_IssueQueueComponent_l187_2 = wokeUpSrc2Mask[2];
  assign when_IssueQueueComponent_l186_3 = wokeUpSrc1Mask[3];
  assign when_IssueQueueComponent_l187_3 = wokeUpSrc2Mask[3];
  assign _zz_1 = ({3'd0,1'b1} <<< issueIdx);
  assign io_allocateIn_fire = (io_allocateIn_valid && io_allocateIn_ready);
  assign _zz_2 = ({3'd0,1'b1} <<< allocateIdx);
  assign _zz_3 = _zz_2[0];
  assign _zz_4 = _zz_2[1];
  assign _zz_5 = _zz_2[2];
  assign _zz_6 = _zz_2[3];
  assign _zz_entriesNext_0_src1Ready = (! io_allocateIn_payload_uop_decoded_useArchSrc1);
  assign _zz_entriesNext_0_src2Ready = (! io_allocateIn_payload_uop_decoded_useArchSrc2);
  assign _zz_7 = ({3'd0,1'b1} <<< allocateIdx);
  assign when_IssueQueueComponent_l212 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l215 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_1 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_1 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_2 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_2 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_3 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_3 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_4 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_4 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_currentValidCount = 3'b000;
  assign _zz_currentValidCount_1 = 3'b001;
  assign _zz_currentValidCount_2 = 3'b001;
  assign _zz_currentValidCount_3 = 3'b010;
  assign _zz_currentValidCount_4 = 3'b001;
  assign _zz_currentValidCount_5 = 3'b010;
  assign _zz_currentValidCount_6 = 3'b010;
  assign _zz_currentValidCount_7 = 3'b011;
  assign currentValidCount = (_zz_currentValidCount_8 + _zz_currentValidCount_10);
  assign logCondition = (io_allocateIn_fire || io_issueOut_fire);
  assign when_IssueQueueComponent_l256 = (logCondition && (3'b000 < currentValidCount));
  always @(posedge clk) begin
    if(reset) begin
      entryValids_0 <= 1'b0;
      entryValids_1 <= 1'b0;
      entryValids_2 <= 1'b0;
      entryValids_3 <= 1'b0;
    end else begin
      entryValids_0 <= entryValidsNext_0;
      entryValids_1 <= entryValidsNext_1;
      entryValids_2 <= entryValidsNext_2;
      entryValids_3 <= entryValidsNext_3;
      if(logCondition) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // IssueQueueComponent.scala:L247
          `else
            if(!1'b0) begin
              $display("NOTE(IssueQueueComponent.scala:247):  [normal] MulEU_IQ-1: STATUS - ValidCount=%x, allocateIn(valid=%x, ready=%x), issueOut(valid=%x, ready=%x)", currentValidCount, io_allocateIn_valid, io_allocateIn_ready, io_issueOut_valid, io_issueOut_ready); // IssueQueueComponent.scala:L247
            end
          `endif
        `endif
      end
      if(when_IssueQueueComponent_l256) begin
        if(entryValids_0) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] MulEU_IQ-1: (LAST CYCLE) ENTRY[0] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_0_robPtr, entries_0_physDest_idx, entries_0_useSrc1, entries_0_src1Tag, entries_0_src1Ready, entries_0_useSrc2, entries_0_src2Tag, entries_0_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_1) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] MulEU_IQ-1: (LAST CYCLE) ENTRY[1] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_1_robPtr, entries_1_physDest_idx, entries_1_useSrc1, entries_1_src1Tag, entries_1_src1Ready, entries_1_useSrc2, entries_1_src2Tag, entries_1_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_2) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] MulEU_IQ-1: (LAST CYCLE) ENTRY[2] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_2_robPtr, entries_2_physDest_idx, entries_2_useSrc1, entries_2_src1Tag, entries_2_src1Ready, entries_2_useSrc2, entries_2_src2Tag, entries_2_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_3) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] MulEU_IQ-1: (LAST CYCLE) ENTRY[3] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_3_robPtr, entries_3_physDest_idx, entries_3_useSrc1, entries_3_src1Tag, entries_3_src1Ready, entries_3_useSrc2, entries_3_src2Tag, entries_3_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
      end
    end
  end

  always @(posedge clk) begin
    entries_0_uop_decoded_pc <= entriesNext_0_uop_decoded_pc;
    entries_0_uop_decoded_isValid <= entriesNext_0_uop_decoded_isValid;
    entries_0_uop_decoded_uopCode <= entriesNext_0_uop_decoded_uopCode;
    entries_0_uop_decoded_exeUnit <= entriesNext_0_uop_decoded_exeUnit;
    entries_0_uop_decoded_isa <= entriesNext_0_uop_decoded_isa;
    entries_0_uop_decoded_archDest_idx <= entriesNext_0_uop_decoded_archDest_idx;
    entries_0_uop_decoded_archDest_rtype <= entriesNext_0_uop_decoded_archDest_rtype;
    entries_0_uop_decoded_writeArchDestEn <= entriesNext_0_uop_decoded_writeArchDestEn;
    entries_0_uop_decoded_archSrc1_idx <= entriesNext_0_uop_decoded_archSrc1_idx;
    entries_0_uop_decoded_archSrc1_rtype <= entriesNext_0_uop_decoded_archSrc1_rtype;
    entries_0_uop_decoded_useArchSrc1 <= entriesNext_0_uop_decoded_useArchSrc1;
    entries_0_uop_decoded_archSrc2_idx <= entriesNext_0_uop_decoded_archSrc2_idx;
    entries_0_uop_decoded_archSrc2_rtype <= entriesNext_0_uop_decoded_archSrc2_rtype;
    entries_0_uop_decoded_useArchSrc2 <= entriesNext_0_uop_decoded_useArchSrc2;
    entries_0_uop_decoded_usePcForAddr <= entriesNext_0_uop_decoded_usePcForAddr;
    entries_0_uop_decoded_imm <= entriesNext_0_uop_decoded_imm;
    entries_0_uop_decoded_immUsage <= entriesNext_0_uop_decoded_immUsage;
    entries_0_uop_decoded_aluCtrl_valid <= entriesNext_0_uop_decoded_aluCtrl_valid;
    entries_0_uop_decoded_aluCtrl_isSub <= entriesNext_0_uop_decoded_aluCtrl_isSub;
    entries_0_uop_decoded_aluCtrl_isAdd <= entriesNext_0_uop_decoded_aluCtrl_isAdd;
    entries_0_uop_decoded_aluCtrl_isSigned <= entriesNext_0_uop_decoded_aluCtrl_isSigned;
    entries_0_uop_decoded_aluCtrl_logicOp <= entriesNext_0_uop_decoded_aluCtrl_logicOp;
    entries_0_uop_decoded_shiftCtrl_valid <= entriesNext_0_uop_decoded_shiftCtrl_valid;
    entries_0_uop_decoded_shiftCtrl_isRight <= entriesNext_0_uop_decoded_shiftCtrl_isRight;
    entries_0_uop_decoded_shiftCtrl_isArithmetic <= entriesNext_0_uop_decoded_shiftCtrl_isArithmetic;
    entries_0_uop_decoded_shiftCtrl_isRotate <= entriesNext_0_uop_decoded_shiftCtrl_isRotate;
    entries_0_uop_decoded_shiftCtrl_isDoubleWord <= entriesNext_0_uop_decoded_shiftCtrl_isDoubleWord;
    entries_0_uop_decoded_mulDivCtrl_valid <= entriesNext_0_uop_decoded_mulDivCtrl_valid;
    entries_0_uop_decoded_mulDivCtrl_isDiv <= entriesNext_0_uop_decoded_mulDivCtrl_isDiv;
    entries_0_uop_decoded_mulDivCtrl_isSigned <= entriesNext_0_uop_decoded_mulDivCtrl_isSigned;
    entries_0_uop_decoded_mulDivCtrl_isWordOp <= entriesNext_0_uop_decoded_mulDivCtrl_isWordOp;
    entries_0_uop_decoded_memCtrl_size <= entriesNext_0_uop_decoded_memCtrl_size;
    entries_0_uop_decoded_memCtrl_isSignedLoad <= entriesNext_0_uop_decoded_memCtrl_isSignedLoad;
    entries_0_uop_decoded_memCtrl_isStore <= entriesNext_0_uop_decoded_memCtrl_isStore;
    entries_0_uop_decoded_memCtrl_isLoadLinked <= entriesNext_0_uop_decoded_memCtrl_isLoadLinked;
    entries_0_uop_decoded_memCtrl_isStoreCond <= entriesNext_0_uop_decoded_memCtrl_isStoreCond;
    entries_0_uop_decoded_memCtrl_atomicOp <= entriesNext_0_uop_decoded_memCtrl_atomicOp;
    entries_0_uop_decoded_memCtrl_isFence <= entriesNext_0_uop_decoded_memCtrl_isFence;
    entries_0_uop_decoded_memCtrl_fenceMode <= entriesNext_0_uop_decoded_memCtrl_fenceMode;
    entries_0_uop_decoded_memCtrl_isCacheOp <= entriesNext_0_uop_decoded_memCtrl_isCacheOp;
    entries_0_uop_decoded_memCtrl_cacheOpType <= entriesNext_0_uop_decoded_memCtrl_cacheOpType;
    entries_0_uop_decoded_memCtrl_isPrefetch <= entriesNext_0_uop_decoded_memCtrl_isPrefetch;
    entries_0_uop_decoded_branchCtrl_condition <= entriesNext_0_uop_decoded_branchCtrl_condition;
    entries_0_uop_decoded_branchCtrl_isJump <= entriesNext_0_uop_decoded_branchCtrl_isJump;
    entries_0_uop_decoded_branchCtrl_isLink <= entriesNext_0_uop_decoded_branchCtrl_isLink;
    entries_0_uop_decoded_branchCtrl_linkReg_idx <= entriesNext_0_uop_decoded_branchCtrl_linkReg_idx;
    entries_0_uop_decoded_branchCtrl_linkReg_rtype <= entriesNext_0_uop_decoded_branchCtrl_linkReg_rtype;
    entries_0_uop_decoded_branchCtrl_isIndirect <= entriesNext_0_uop_decoded_branchCtrl_isIndirect;
    entries_0_uop_decoded_branchCtrl_laCfIdx <= entriesNext_0_uop_decoded_branchCtrl_laCfIdx;
    entries_0_uop_decoded_fpuCtrl_opType <= entriesNext_0_uop_decoded_fpuCtrl_opType;
    entries_0_uop_decoded_fpuCtrl_fpSizeSrc1 <= entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc1;
    entries_0_uop_decoded_fpuCtrl_fpSizeSrc2 <= entriesNext_0_uop_decoded_fpuCtrl_fpSizeSrc2;
    entries_0_uop_decoded_fpuCtrl_fpSizeDest <= entriesNext_0_uop_decoded_fpuCtrl_fpSizeDest;
    entries_0_uop_decoded_fpuCtrl_roundingMode <= entriesNext_0_uop_decoded_fpuCtrl_roundingMode;
    entries_0_uop_decoded_fpuCtrl_isIntegerDest <= entriesNext_0_uop_decoded_fpuCtrl_isIntegerDest;
    entries_0_uop_decoded_fpuCtrl_isSignedCvt <= entriesNext_0_uop_decoded_fpuCtrl_isSignedCvt;
    entries_0_uop_decoded_fpuCtrl_fmaNegSrc1 <= entriesNext_0_uop_decoded_fpuCtrl_fmaNegSrc1;
    entries_0_uop_decoded_fpuCtrl_fcmpCond <= entriesNext_0_uop_decoded_fpuCtrl_fcmpCond;
    entries_0_uop_decoded_csrCtrl_csrAddr <= entriesNext_0_uop_decoded_csrCtrl_csrAddr;
    entries_0_uop_decoded_csrCtrl_isWrite <= entriesNext_0_uop_decoded_csrCtrl_isWrite;
    entries_0_uop_decoded_csrCtrl_isRead <= entriesNext_0_uop_decoded_csrCtrl_isRead;
    entries_0_uop_decoded_csrCtrl_isExchange <= entriesNext_0_uop_decoded_csrCtrl_isExchange;
    entries_0_uop_decoded_csrCtrl_useUimmAsSrc <= entriesNext_0_uop_decoded_csrCtrl_useUimmAsSrc;
    entries_0_uop_decoded_sysCtrl_sysCode <= entriesNext_0_uop_decoded_sysCtrl_sysCode;
    entries_0_uop_decoded_sysCtrl_isExceptionReturn <= entriesNext_0_uop_decoded_sysCtrl_isExceptionReturn;
    entries_0_uop_decoded_sysCtrl_isTlbOp <= entriesNext_0_uop_decoded_sysCtrl_isTlbOp;
    entries_0_uop_decoded_sysCtrl_tlbOpType <= entriesNext_0_uop_decoded_sysCtrl_tlbOpType;
    entries_0_uop_decoded_decodeExceptionCode <= entriesNext_0_uop_decoded_decodeExceptionCode;
    entries_0_uop_decoded_hasDecodeException <= entriesNext_0_uop_decoded_hasDecodeException;
    entries_0_uop_decoded_isMicrocode <= entriesNext_0_uop_decoded_isMicrocode;
    entries_0_uop_decoded_microcodeEntry <= entriesNext_0_uop_decoded_microcodeEntry;
    entries_0_uop_decoded_isSerializing <= entriesNext_0_uop_decoded_isSerializing;
    entries_0_uop_decoded_isBranchOrJump <= entriesNext_0_uop_decoded_isBranchOrJump;
    entries_0_uop_decoded_branchPrediction_isTaken <= entriesNext_0_uop_decoded_branchPrediction_isTaken;
    entries_0_uop_decoded_branchPrediction_target <= entriesNext_0_uop_decoded_branchPrediction_target;
    entries_0_uop_decoded_branchPrediction_wasPredicted <= entriesNext_0_uop_decoded_branchPrediction_wasPredicted;
    entries_0_uop_rename_physSrc1_idx <= entriesNext_0_uop_rename_physSrc1_idx;
    entries_0_uop_rename_physSrc1IsFpr <= entriesNext_0_uop_rename_physSrc1IsFpr;
    entries_0_uop_rename_physSrc2_idx <= entriesNext_0_uop_rename_physSrc2_idx;
    entries_0_uop_rename_physSrc2IsFpr <= entriesNext_0_uop_rename_physSrc2IsFpr;
    entries_0_uop_rename_physDest_idx <= entriesNext_0_uop_rename_physDest_idx;
    entries_0_uop_rename_physDestIsFpr <= entriesNext_0_uop_rename_physDestIsFpr;
    entries_0_uop_rename_oldPhysDest_idx <= entriesNext_0_uop_rename_oldPhysDest_idx;
    entries_0_uop_rename_oldPhysDestIsFpr <= entriesNext_0_uop_rename_oldPhysDestIsFpr;
    entries_0_uop_rename_allocatesPhysDest <= entriesNext_0_uop_rename_allocatesPhysDest;
    entries_0_uop_rename_writesToPhysReg <= entriesNext_0_uop_rename_writesToPhysReg;
    entries_0_uop_robPtr <= entriesNext_0_uop_robPtr;
    entries_0_uop_uniqueId <= entriesNext_0_uop_uniqueId;
    entries_0_uop_dispatched <= entriesNext_0_uop_dispatched;
    entries_0_uop_executed <= entriesNext_0_uop_executed;
    entries_0_uop_hasException <= entriesNext_0_uop_hasException;
    entries_0_uop_exceptionCode <= entriesNext_0_uop_exceptionCode;
    entries_0_robPtr <= entriesNext_0_robPtr;
    entries_0_physDest_idx <= entriesNext_0_physDest_idx;
    entries_0_physDestIsFpr <= entriesNext_0_physDestIsFpr;
    entries_0_writesToPhysReg <= entriesNext_0_writesToPhysReg;
    entries_0_useSrc1 <= entriesNext_0_useSrc1;
    entries_0_src1Data <= entriesNext_0_src1Data;
    entries_0_src1Tag <= entriesNext_0_src1Tag;
    entries_0_src1Ready <= entriesNext_0_src1Ready;
    entries_0_src1IsFpr <= entriesNext_0_src1IsFpr;
    entries_0_useSrc2 <= entriesNext_0_useSrc2;
    entries_0_src2Data <= entriesNext_0_src2Data;
    entries_0_src2Tag <= entriesNext_0_src2Tag;
    entries_0_src2Ready <= entriesNext_0_src2Ready;
    entries_0_src2IsFpr <= entriesNext_0_src2IsFpr;
    entries_0_mulDivCtrl_valid <= entriesNext_0_mulDivCtrl_valid;
    entries_0_mulDivCtrl_isDiv <= entriesNext_0_mulDivCtrl_isDiv;
    entries_0_mulDivCtrl_isSigned <= entriesNext_0_mulDivCtrl_isSigned;
    entries_0_mulDivCtrl_isWordOp <= entriesNext_0_mulDivCtrl_isWordOp;
    entries_1_uop_decoded_pc <= entriesNext_1_uop_decoded_pc;
    entries_1_uop_decoded_isValid <= entriesNext_1_uop_decoded_isValid;
    entries_1_uop_decoded_uopCode <= entriesNext_1_uop_decoded_uopCode;
    entries_1_uop_decoded_exeUnit <= entriesNext_1_uop_decoded_exeUnit;
    entries_1_uop_decoded_isa <= entriesNext_1_uop_decoded_isa;
    entries_1_uop_decoded_archDest_idx <= entriesNext_1_uop_decoded_archDest_idx;
    entries_1_uop_decoded_archDest_rtype <= entriesNext_1_uop_decoded_archDest_rtype;
    entries_1_uop_decoded_writeArchDestEn <= entriesNext_1_uop_decoded_writeArchDestEn;
    entries_1_uop_decoded_archSrc1_idx <= entriesNext_1_uop_decoded_archSrc1_idx;
    entries_1_uop_decoded_archSrc1_rtype <= entriesNext_1_uop_decoded_archSrc1_rtype;
    entries_1_uop_decoded_useArchSrc1 <= entriesNext_1_uop_decoded_useArchSrc1;
    entries_1_uop_decoded_archSrc2_idx <= entriesNext_1_uop_decoded_archSrc2_idx;
    entries_1_uop_decoded_archSrc2_rtype <= entriesNext_1_uop_decoded_archSrc2_rtype;
    entries_1_uop_decoded_useArchSrc2 <= entriesNext_1_uop_decoded_useArchSrc2;
    entries_1_uop_decoded_usePcForAddr <= entriesNext_1_uop_decoded_usePcForAddr;
    entries_1_uop_decoded_imm <= entriesNext_1_uop_decoded_imm;
    entries_1_uop_decoded_immUsage <= entriesNext_1_uop_decoded_immUsage;
    entries_1_uop_decoded_aluCtrl_valid <= entriesNext_1_uop_decoded_aluCtrl_valid;
    entries_1_uop_decoded_aluCtrl_isSub <= entriesNext_1_uop_decoded_aluCtrl_isSub;
    entries_1_uop_decoded_aluCtrl_isAdd <= entriesNext_1_uop_decoded_aluCtrl_isAdd;
    entries_1_uop_decoded_aluCtrl_isSigned <= entriesNext_1_uop_decoded_aluCtrl_isSigned;
    entries_1_uop_decoded_aluCtrl_logicOp <= entriesNext_1_uop_decoded_aluCtrl_logicOp;
    entries_1_uop_decoded_shiftCtrl_valid <= entriesNext_1_uop_decoded_shiftCtrl_valid;
    entries_1_uop_decoded_shiftCtrl_isRight <= entriesNext_1_uop_decoded_shiftCtrl_isRight;
    entries_1_uop_decoded_shiftCtrl_isArithmetic <= entriesNext_1_uop_decoded_shiftCtrl_isArithmetic;
    entries_1_uop_decoded_shiftCtrl_isRotate <= entriesNext_1_uop_decoded_shiftCtrl_isRotate;
    entries_1_uop_decoded_shiftCtrl_isDoubleWord <= entriesNext_1_uop_decoded_shiftCtrl_isDoubleWord;
    entries_1_uop_decoded_mulDivCtrl_valid <= entriesNext_1_uop_decoded_mulDivCtrl_valid;
    entries_1_uop_decoded_mulDivCtrl_isDiv <= entriesNext_1_uop_decoded_mulDivCtrl_isDiv;
    entries_1_uop_decoded_mulDivCtrl_isSigned <= entriesNext_1_uop_decoded_mulDivCtrl_isSigned;
    entries_1_uop_decoded_mulDivCtrl_isWordOp <= entriesNext_1_uop_decoded_mulDivCtrl_isWordOp;
    entries_1_uop_decoded_memCtrl_size <= entriesNext_1_uop_decoded_memCtrl_size;
    entries_1_uop_decoded_memCtrl_isSignedLoad <= entriesNext_1_uop_decoded_memCtrl_isSignedLoad;
    entries_1_uop_decoded_memCtrl_isStore <= entriesNext_1_uop_decoded_memCtrl_isStore;
    entries_1_uop_decoded_memCtrl_isLoadLinked <= entriesNext_1_uop_decoded_memCtrl_isLoadLinked;
    entries_1_uop_decoded_memCtrl_isStoreCond <= entriesNext_1_uop_decoded_memCtrl_isStoreCond;
    entries_1_uop_decoded_memCtrl_atomicOp <= entriesNext_1_uop_decoded_memCtrl_atomicOp;
    entries_1_uop_decoded_memCtrl_isFence <= entriesNext_1_uop_decoded_memCtrl_isFence;
    entries_1_uop_decoded_memCtrl_fenceMode <= entriesNext_1_uop_decoded_memCtrl_fenceMode;
    entries_1_uop_decoded_memCtrl_isCacheOp <= entriesNext_1_uop_decoded_memCtrl_isCacheOp;
    entries_1_uop_decoded_memCtrl_cacheOpType <= entriesNext_1_uop_decoded_memCtrl_cacheOpType;
    entries_1_uop_decoded_memCtrl_isPrefetch <= entriesNext_1_uop_decoded_memCtrl_isPrefetch;
    entries_1_uop_decoded_branchCtrl_condition <= entriesNext_1_uop_decoded_branchCtrl_condition;
    entries_1_uop_decoded_branchCtrl_isJump <= entriesNext_1_uop_decoded_branchCtrl_isJump;
    entries_1_uop_decoded_branchCtrl_isLink <= entriesNext_1_uop_decoded_branchCtrl_isLink;
    entries_1_uop_decoded_branchCtrl_linkReg_idx <= entriesNext_1_uop_decoded_branchCtrl_linkReg_idx;
    entries_1_uop_decoded_branchCtrl_linkReg_rtype <= entriesNext_1_uop_decoded_branchCtrl_linkReg_rtype;
    entries_1_uop_decoded_branchCtrl_isIndirect <= entriesNext_1_uop_decoded_branchCtrl_isIndirect;
    entries_1_uop_decoded_branchCtrl_laCfIdx <= entriesNext_1_uop_decoded_branchCtrl_laCfIdx;
    entries_1_uop_decoded_fpuCtrl_opType <= entriesNext_1_uop_decoded_fpuCtrl_opType;
    entries_1_uop_decoded_fpuCtrl_fpSizeSrc1 <= entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc1;
    entries_1_uop_decoded_fpuCtrl_fpSizeSrc2 <= entriesNext_1_uop_decoded_fpuCtrl_fpSizeSrc2;
    entries_1_uop_decoded_fpuCtrl_fpSizeDest <= entriesNext_1_uop_decoded_fpuCtrl_fpSizeDest;
    entries_1_uop_decoded_fpuCtrl_roundingMode <= entriesNext_1_uop_decoded_fpuCtrl_roundingMode;
    entries_1_uop_decoded_fpuCtrl_isIntegerDest <= entriesNext_1_uop_decoded_fpuCtrl_isIntegerDest;
    entries_1_uop_decoded_fpuCtrl_isSignedCvt <= entriesNext_1_uop_decoded_fpuCtrl_isSignedCvt;
    entries_1_uop_decoded_fpuCtrl_fmaNegSrc1 <= entriesNext_1_uop_decoded_fpuCtrl_fmaNegSrc1;
    entries_1_uop_decoded_fpuCtrl_fcmpCond <= entriesNext_1_uop_decoded_fpuCtrl_fcmpCond;
    entries_1_uop_decoded_csrCtrl_csrAddr <= entriesNext_1_uop_decoded_csrCtrl_csrAddr;
    entries_1_uop_decoded_csrCtrl_isWrite <= entriesNext_1_uop_decoded_csrCtrl_isWrite;
    entries_1_uop_decoded_csrCtrl_isRead <= entriesNext_1_uop_decoded_csrCtrl_isRead;
    entries_1_uop_decoded_csrCtrl_isExchange <= entriesNext_1_uop_decoded_csrCtrl_isExchange;
    entries_1_uop_decoded_csrCtrl_useUimmAsSrc <= entriesNext_1_uop_decoded_csrCtrl_useUimmAsSrc;
    entries_1_uop_decoded_sysCtrl_sysCode <= entriesNext_1_uop_decoded_sysCtrl_sysCode;
    entries_1_uop_decoded_sysCtrl_isExceptionReturn <= entriesNext_1_uop_decoded_sysCtrl_isExceptionReturn;
    entries_1_uop_decoded_sysCtrl_isTlbOp <= entriesNext_1_uop_decoded_sysCtrl_isTlbOp;
    entries_1_uop_decoded_sysCtrl_tlbOpType <= entriesNext_1_uop_decoded_sysCtrl_tlbOpType;
    entries_1_uop_decoded_decodeExceptionCode <= entriesNext_1_uop_decoded_decodeExceptionCode;
    entries_1_uop_decoded_hasDecodeException <= entriesNext_1_uop_decoded_hasDecodeException;
    entries_1_uop_decoded_isMicrocode <= entriesNext_1_uop_decoded_isMicrocode;
    entries_1_uop_decoded_microcodeEntry <= entriesNext_1_uop_decoded_microcodeEntry;
    entries_1_uop_decoded_isSerializing <= entriesNext_1_uop_decoded_isSerializing;
    entries_1_uop_decoded_isBranchOrJump <= entriesNext_1_uop_decoded_isBranchOrJump;
    entries_1_uop_decoded_branchPrediction_isTaken <= entriesNext_1_uop_decoded_branchPrediction_isTaken;
    entries_1_uop_decoded_branchPrediction_target <= entriesNext_1_uop_decoded_branchPrediction_target;
    entries_1_uop_decoded_branchPrediction_wasPredicted <= entriesNext_1_uop_decoded_branchPrediction_wasPredicted;
    entries_1_uop_rename_physSrc1_idx <= entriesNext_1_uop_rename_physSrc1_idx;
    entries_1_uop_rename_physSrc1IsFpr <= entriesNext_1_uop_rename_physSrc1IsFpr;
    entries_1_uop_rename_physSrc2_idx <= entriesNext_1_uop_rename_physSrc2_idx;
    entries_1_uop_rename_physSrc2IsFpr <= entriesNext_1_uop_rename_physSrc2IsFpr;
    entries_1_uop_rename_physDest_idx <= entriesNext_1_uop_rename_physDest_idx;
    entries_1_uop_rename_physDestIsFpr <= entriesNext_1_uop_rename_physDestIsFpr;
    entries_1_uop_rename_oldPhysDest_idx <= entriesNext_1_uop_rename_oldPhysDest_idx;
    entries_1_uop_rename_oldPhysDestIsFpr <= entriesNext_1_uop_rename_oldPhysDestIsFpr;
    entries_1_uop_rename_allocatesPhysDest <= entriesNext_1_uop_rename_allocatesPhysDest;
    entries_1_uop_rename_writesToPhysReg <= entriesNext_1_uop_rename_writesToPhysReg;
    entries_1_uop_robPtr <= entriesNext_1_uop_robPtr;
    entries_1_uop_uniqueId <= entriesNext_1_uop_uniqueId;
    entries_1_uop_dispatched <= entriesNext_1_uop_dispatched;
    entries_1_uop_executed <= entriesNext_1_uop_executed;
    entries_1_uop_hasException <= entriesNext_1_uop_hasException;
    entries_1_uop_exceptionCode <= entriesNext_1_uop_exceptionCode;
    entries_1_robPtr <= entriesNext_1_robPtr;
    entries_1_physDest_idx <= entriesNext_1_physDest_idx;
    entries_1_physDestIsFpr <= entriesNext_1_physDestIsFpr;
    entries_1_writesToPhysReg <= entriesNext_1_writesToPhysReg;
    entries_1_useSrc1 <= entriesNext_1_useSrc1;
    entries_1_src1Data <= entriesNext_1_src1Data;
    entries_1_src1Tag <= entriesNext_1_src1Tag;
    entries_1_src1Ready <= entriesNext_1_src1Ready;
    entries_1_src1IsFpr <= entriesNext_1_src1IsFpr;
    entries_1_useSrc2 <= entriesNext_1_useSrc2;
    entries_1_src2Data <= entriesNext_1_src2Data;
    entries_1_src2Tag <= entriesNext_1_src2Tag;
    entries_1_src2Ready <= entriesNext_1_src2Ready;
    entries_1_src2IsFpr <= entriesNext_1_src2IsFpr;
    entries_1_mulDivCtrl_valid <= entriesNext_1_mulDivCtrl_valid;
    entries_1_mulDivCtrl_isDiv <= entriesNext_1_mulDivCtrl_isDiv;
    entries_1_mulDivCtrl_isSigned <= entriesNext_1_mulDivCtrl_isSigned;
    entries_1_mulDivCtrl_isWordOp <= entriesNext_1_mulDivCtrl_isWordOp;
    entries_2_uop_decoded_pc <= entriesNext_2_uop_decoded_pc;
    entries_2_uop_decoded_isValid <= entriesNext_2_uop_decoded_isValid;
    entries_2_uop_decoded_uopCode <= entriesNext_2_uop_decoded_uopCode;
    entries_2_uop_decoded_exeUnit <= entriesNext_2_uop_decoded_exeUnit;
    entries_2_uop_decoded_isa <= entriesNext_2_uop_decoded_isa;
    entries_2_uop_decoded_archDest_idx <= entriesNext_2_uop_decoded_archDest_idx;
    entries_2_uop_decoded_archDest_rtype <= entriesNext_2_uop_decoded_archDest_rtype;
    entries_2_uop_decoded_writeArchDestEn <= entriesNext_2_uop_decoded_writeArchDestEn;
    entries_2_uop_decoded_archSrc1_idx <= entriesNext_2_uop_decoded_archSrc1_idx;
    entries_2_uop_decoded_archSrc1_rtype <= entriesNext_2_uop_decoded_archSrc1_rtype;
    entries_2_uop_decoded_useArchSrc1 <= entriesNext_2_uop_decoded_useArchSrc1;
    entries_2_uop_decoded_archSrc2_idx <= entriesNext_2_uop_decoded_archSrc2_idx;
    entries_2_uop_decoded_archSrc2_rtype <= entriesNext_2_uop_decoded_archSrc2_rtype;
    entries_2_uop_decoded_useArchSrc2 <= entriesNext_2_uop_decoded_useArchSrc2;
    entries_2_uop_decoded_usePcForAddr <= entriesNext_2_uop_decoded_usePcForAddr;
    entries_2_uop_decoded_imm <= entriesNext_2_uop_decoded_imm;
    entries_2_uop_decoded_immUsage <= entriesNext_2_uop_decoded_immUsage;
    entries_2_uop_decoded_aluCtrl_valid <= entriesNext_2_uop_decoded_aluCtrl_valid;
    entries_2_uop_decoded_aluCtrl_isSub <= entriesNext_2_uop_decoded_aluCtrl_isSub;
    entries_2_uop_decoded_aluCtrl_isAdd <= entriesNext_2_uop_decoded_aluCtrl_isAdd;
    entries_2_uop_decoded_aluCtrl_isSigned <= entriesNext_2_uop_decoded_aluCtrl_isSigned;
    entries_2_uop_decoded_aluCtrl_logicOp <= entriesNext_2_uop_decoded_aluCtrl_logicOp;
    entries_2_uop_decoded_shiftCtrl_valid <= entriesNext_2_uop_decoded_shiftCtrl_valid;
    entries_2_uop_decoded_shiftCtrl_isRight <= entriesNext_2_uop_decoded_shiftCtrl_isRight;
    entries_2_uop_decoded_shiftCtrl_isArithmetic <= entriesNext_2_uop_decoded_shiftCtrl_isArithmetic;
    entries_2_uop_decoded_shiftCtrl_isRotate <= entriesNext_2_uop_decoded_shiftCtrl_isRotate;
    entries_2_uop_decoded_shiftCtrl_isDoubleWord <= entriesNext_2_uop_decoded_shiftCtrl_isDoubleWord;
    entries_2_uop_decoded_mulDivCtrl_valid <= entriesNext_2_uop_decoded_mulDivCtrl_valid;
    entries_2_uop_decoded_mulDivCtrl_isDiv <= entriesNext_2_uop_decoded_mulDivCtrl_isDiv;
    entries_2_uop_decoded_mulDivCtrl_isSigned <= entriesNext_2_uop_decoded_mulDivCtrl_isSigned;
    entries_2_uop_decoded_mulDivCtrl_isWordOp <= entriesNext_2_uop_decoded_mulDivCtrl_isWordOp;
    entries_2_uop_decoded_memCtrl_size <= entriesNext_2_uop_decoded_memCtrl_size;
    entries_2_uop_decoded_memCtrl_isSignedLoad <= entriesNext_2_uop_decoded_memCtrl_isSignedLoad;
    entries_2_uop_decoded_memCtrl_isStore <= entriesNext_2_uop_decoded_memCtrl_isStore;
    entries_2_uop_decoded_memCtrl_isLoadLinked <= entriesNext_2_uop_decoded_memCtrl_isLoadLinked;
    entries_2_uop_decoded_memCtrl_isStoreCond <= entriesNext_2_uop_decoded_memCtrl_isStoreCond;
    entries_2_uop_decoded_memCtrl_atomicOp <= entriesNext_2_uop_decoded_memCtrl_atomicOp;
    entries_2_uop_decoded_memCtrl_isFence <= entriesNext_2_uop_decoded_memCtrl_isFence;
    entries_2_uop_decoded_memCtrl_fenceMode <= entriesNext_2_uop_decoded_memCtrl_fenceMode;
    entries_2_uop_decoded_memCtrl_isCacheOp <= entriesNext_2_uop_decoded_memCtrl_isCacheOp;
    entries_2_uop_decoded_memCtrl_cacheOpType <= entriesNext_2_uop_decoded_memCtrl_cacheOpType;
    entries_2_uop_decoded_memCtrl_isPrefetch <= entriesNext_2_uop_decoded_memCtrl_isPrefetch;
    entries_2_uop_decoded_branchCtrl_condition <= entriesNext_2_uop_decoded_branchCtrl_condition;
    entries_2_uop_decoded_branchCtrl_isJump <= entriesNext_2_uop_decoded_branchCtrl_isJump;
    entries_2_uop_decoded_branchCtrl_isLink <= entriesNext_2_uop_decoded_branchCtrl_isLink;
    entries_2_uop_decoded_branchCtrl_linkReg_idx <= entriesNext_2_uop_decoded_branchCtrl_linkReg_idx;
    entries_2_uop_decoded_branchCtrl_linkReg_rtype <= entriesNext_2_uop_decoded_branchCtrl_linkReg_rtype;
    entries_2_uop_decoded_branchCtrl_isIndirect <= entriesNext_2_uop_decoded_branchCtrl_isIndirect;
    entries_2_uop_decoded_branchCtrl_laCfIdx <= entriesNext_2_uop_decoded_branchCtrl_laCfIdx;
    entries_2_uop_decoded_fpuCtrl_opType <= entriesNext_2_uop_decoded_fpuCtrl_opType;
    entries_2_uop_decoded_fpuCtrl_fpSizeSrc1 <= entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc1;
    entries_2_uop_decoded_fpuCtrl_fpSizeSrc2 <= entriesNext_2_uop_decoded_fpuCtrl_fpSizeSrc2;
    entries_2_uop_decoded_fpuCtrl_fpSizeDest <= entriesNext_2_uop_decoded_fpuCtrl_fpSizeDest;
    entries_2_uop_decoded_fpuCtrl_roundingMode <= entriesNext_2_uop_decoded_fpuCtrl_roundingMode;
    entries_2_uop_decoded_fpuCtrl_isIntegerDest <= entriesNext_2_uop_decoded_fpuCtrl_isIntegerDest;
    entries_2_uop_decoded_fpuCtrl_isSignedCvt <= entriesNext_2_uop_decoded_fpuCtrl_isSignedCvt;
    entries_2_uop_decoded_fpuCtrl_fmaNegSrc1 <= entriesNext_2_uop_decoded_fpuCtrl_fmaNegSrc1;
    entries_2_uop_decoded_fpuCtrl_fcmpCond <= entriesNext_2_uop_decoded_fpuCtrl_fcmpCond;
    entries_2_uop_decoded_csrCtrl_csrAddr <= entriesNext_2_uop_decoded_csrCtrl_csrAddr;
    entries_2_uop_decoded_csrCtrl_isWrite <= entriesNext_2_uop_decoded_csrCtrl_isWrite;
    entries_2_uop_decoded_csrCtrl_isRead <= entriesNext_2_uop_decoded_csrCtrl_isRead;
    entries_2_uop_decoded_csrCtrl_isExchange <= entriesNext_2_uop_decoded_csrCtrl_isExchange;
    entries_2_uop_decoded_csrCtrl_useUimmAsSrc <= entriesNext_2_uop_decoded_csrCtrl_useUimmAsSrc;
    entries_2_uop_decoded_sysCtrl_sysCode <= entriesNext_2_uop_decoded_sysCtrl_sysCode;
    entries_2_uop_decoded_sysCtrl_isExceptionReturn <= entriesNext_2_uop_decoded_sysCtrl_isExceptionReturn;
    entries_2_uop_decoded_sysCtrl_isTlbOp <= entriesNext_2_uop_decoded_sysCtrl_isTlbOp;
    entries_2_uop_decoded_sysCtrl_tlbOpType <= entriesNext_2_uop_decoded_sysCtrl_tlbOpType;
    entries_2_uop_decoded_decodeExceptionCode <= entriesNext_2_uop_decoded_decodeExceptionCode;
    entries_2_uop_decoded_hasDecodeException <= entriesNext_2_uop_decoded_hasDecodeException;
    entries_2_uop_decoded_isMicrocode <= entriesNext_2_uop_decoded_isMicrocode;
    entries_2_uop_decoded_microcodeEntry <= entriesNext_2_uop_decoded_microcodeEntry;
    entries_2_uop_decoded_isSerializing <= entriesNext_2_uop_decoded_isSerializing;
    entries_2_uop_decoded_isBranchOrJump <= entriesNext_2_uop_decoded_isBranchOrJump;
    entries_2_uop_decoded_branchPrediction_isTaken <= entriesNext_2_uop_decoded_branchPrediction_isTaken;
    entries_2_uop_decoded_branchPrediction_target <= entriesNext_2_uop_decoded_branchPrediction_target;
    entries_2_uop_decoded_branchPrediction_wasPredicted <= entriesNext_2_uop_decoded_branchPrediction_wasPredicted;
    entries_2_uop_rename_physSrc1_idx <= entriesNext_2_uop_rename_physSrc1_idx;
    entries_2_uop_rename_physSrc1IsFpr <= entriesNext_2_uop_rename_physSrc1IsFpr;
    entries_2_uop_rename_physSrc2_idx <= entriesNext_2_uop_rename_physSrc2_idx;
    entries_2_uop_rename_physSrc2IsFpr <= entriesNext_2_uop_rename_physSrc2IsFpr;
    entries_2_uop_rename_physDest_idx <= entriesNext_2_uop_rename_physDest_idx;
    entries_2_uop_rename_physDestIsFpr <= entriesNext_2_uop_rename_physDestIsFpr;
    entries_2_uop_rename_oldPhysDest_idx <= entriesNext_2_uop_rename_oldPhysDest_idx;
    entries_2_uop_rename_oldPhysDestIsFpr <= entriesNext_2_uop_rename_oldPhysDestIsFpr;
    entries_2_uop_rename_allocatesPhysDest <= entriesNext_2_uop_rename_allocatesPhysDest;
    entries_2_uop_rename_writesToPhysReg <= entriesNext_2_uop_rename_writesToPhysReg;
    entries_2_uop_robPtr <= entriesNext_2_uop_robPtr;
    entries_2_uop_uniqueId <= entriesNext_2_uop_uniqueId;
    entries_2_uop_dispatched <= entriesNext_2_uop_dispatched;
    entries_2_uop_executed <= entriesNext_2_uop_executed;
    entries_2_uop_hasException <= entriesNext_2_uop_hasException;
    entries_2_uop_exceptionCode <= entriesNext_2_uop_exceptionCode;
    entries_2_robPtr <= entriesNext_2_robPtr;
    entries_2_physDest_idx <= entriesNext_2_physDest_idx;
    entries_2_physDestIsFpr <= entriesNext_2_physDestIsFpr;
    entries_2_writesToPhysReg <= entriesNext_2_writesToPhysReg;
    entries_2_useSrc1 <= entriesNext_2_useSrc1;
    entries_2_src1Data <= entriesNext_2_src1Data;
    entries_2_src1Tag <= entriesNext_2_src1Tag;
    entries_2_src1Ready <= entriesNext_2_src1Ready;
    entries_2_src1IsFpr <= entriesNext_2_src1IsFpr;
    entries_2_useSrc2 <= entriesNext_2_useSrc2;
    entries_2_src2Data <= entriesNext_2_src2Data;
    entries_2_src2Tag <= entriesNext_2_src2Tag;
    entries_2_src2Ready <= entriesNext_2_src2Ready;
    entries_2_src2IsFpr <= entriesNext_2_src2IsFpr;
    entries_2_mulDivCtrl_valid <= entriesNext_2_mulDivCtrl_valid;
    entries_2_mulDivCtrl_isDiv <= entriesNext_2_mulDivCtrl_isDiv;
    entries_2_mulDivCtrl_isSigned <= entriesNext_2_mulDivCtrl_isSigned;
    entries_2_mulDivCtrl_isWordOp <= entriesNext_2_mulDivCtrl_isWordOp;
    entries_3_uop_decoded_pc <= entriesNext_3_uop_decoded_pc;
    entries_3_uop_decoded_isValid <= entriesNext_3_uop_decoded_isValid;
    entries_3_uop_decoded_uopCode <= entriesNext_3_uop_decoded_uopCode;
    entries_3_uop_decoded_exeUnit <= entriesNext_3_uop_decoded_exeUnit;
    entries_3_uop_decoded_isa <= entriesNext_3_uop_decoded_isa;
    entries_3_uop_decoded_archDest_idx <= entriesNext_3_uop_decoded_archDest_idx;
    entries_3_uop_decoded_archDest_rtype <= entriesNext_3_uop_decoded_archDest_rtype;
    entries_3_uop_decoded_writeArchDestEn <= entriesNext_3_uop_decoded_writeArchDestEn;
    entries_3_uop_decoded_archSrc1_idx <= entriesNext_3_uop_decoded_archSrc1_idx;
    entries_3_uop_decoded_archSrc1_rtype <= entriesNext_3_uop_decoded_archSrc1_rtype;
    entries_3_uop_decoded_useArchSrc1 <= entriesNext_3_uop_decoded_useArchSrc1;
    entries_3_uop_decoded_archSrc2_idx <= entriesNext_3_uop_decoded_archSrc2_idx;
    entries_3_uop_decoded_archSrc2_rtype <= entriesNext_3_uop_decoded_archSrc2_rtype;
    entries_3_uop_decoded_useArchSrc2 <= entriesNext_3_uop_decoded_useArchSrc2;
    entries_3_uop_decoded_usePcForAddr <= entriesNext_3_uop_decoded_usePcForAddr;
    entries_3_uop_decoded_imm <= entriesNext_3_uop_decoded_imm;
    entries_3_uop_decoded_immUsage <= entriesNext_3_uop_decoded_immUsage;
    entries_3_uop_decoded_aluCtrl_valid <= entriesNext_3_uop_decoded_aluCtrl_valid;
    entries_3_uop_decoded_aluCtrl_isSub <= entriesNext_3_uop_decoded_aluCtrl_isSub;
    entries_3_uop_decoded_aluCtrl_isAdd <= entriesNext_3_uop_decoded_aluCtrl_isAdd;
    entries_3_uop_decoded_aluCtrl_isSigned <= entriesNext_3_uop_decoded_aluCtrl_isSigned;
    entries_3_uop_decoded_aluCtrl_logicOp <= entriesNext_3_uop_decoded_aluCtrl_logicOp;
    entries_3_uop_decoded_shiftCtrl_valid <= entriesNext_3_uop_decoded_shiftCtrl_valid;
    entries_3_uop_decoded_shiftCtrl_isRight <= entriesNext_3_uop_decoded_shiftCtrl_isRight;
    entries_3_uop_decoded_shiftCtrl_isArithmetic <= entriesNext_3_uop_decoded_shiftCtrl_isArithmetic;
    entries_3_uop_decoded_shiftCtrl_isRotate <= entriesNext_3_uop_decoded_shiftCtrl_isRotate;
    entries_3_uop_decoded_shiftCtrl_isDoubleWord <= entriesNext_3_uop_decoded_shiftCtrl_isDoubleWord;
    entries_3_uop_decoded_mulDivCtrl_valid <= entriesNext_3_uop_decoded_mulDivCtrl_valid;
    entries_3_uop_decoded_mulDivCtrl_isDiv <= entriesNext_3_uop_decoded_mulDivCtrl_isDiv;
    entries_3_uop_decoded_mulDivCtrl_isSigned <= entriesNext_3_uop_decoded_mulDivCtrl_isSigned;
    entries_3_uop_decoded_mulDivCtrl_isWordOp <= entriesNext_3_uop_decoded_mulDivCtrl_isWordOp;
    entries_3_uop_decoded_memCtrl_size <= entriesNext_3_uop_decoded_memCtrl_size;
    entries_3_uop_decoded_memCtrl_isSignedLoad <= entriesNext_3_uop_decoded_memCtrl_isSignedLoad;
    entries_3_uop_decoded_memCtrl_isStore <= entriesNext_3_uop_decoded_memCtrl_isStore;
    entries_3_uop_decoded_memCtrl_isLoadLinked <= entriesNext_3_uop_decoded_memCtrl_isLoadLinked;
    entries_3_uop_decoded_memCtrl_isStoreCond <= entriesNext_3_uop_decoded_memCtrl_isStoreCond;
    entries_3_uop_decoded_memCtrl_atomicOp <= entriesNext_3_uop_decoded_memCtrl_atomicOp;
    entries_3_uop_decoded_memCtrl_isFence <= entriesNext_3_uop_decoded_memCtrl_isFence;
    entries_3_uop_decoded_memCtrl_fenceMode <= entriesNext_3_uop_decoded_memCtrl_fenceMode;
    entries_3_uop_decoded_memCtrl_isCacheOp <= entriesNext_3_uop_decoded_memCtrl_isCacheOp;
    entries_3_uop_decoded_memCtrl_cacheOpType <= entriesNext_3_uop_decoded_memCtrl_cacheOpType;
    entries_3_uop_decoded_memCtrl_isPrefetch <= entriesNext_3_uop_decoded_memCtrl_isPrefetch;
    entries_3_uop_decoded_branchCtrl_condition <= entriesNext_3_uop_decoded_branchCtrl_condition;
    entries_3_uop_decoded_branchCtrl_isJump <= entriesNext_3_uop_decoded_branchCtrl_isJump;
    entries_3_uop_decoded_branchCtrl_isLink <= entriesNext_3_uop_decoded_branchCtrl_isLink;
    entries_3_uop_decoded_branchCtrl_linkReg_idx <= entriesNext_3_uop_decoded_branchCtrl_linkReg_idx;
    entries_3_uop_decoded_branchCtrl_linkReg_rtype <= entriesNext_3_uop_decoded_branchCtrl_linkReg_rtype;
    entries_3_uop_decoded_branchCtrl_isIndirect <= entriesNext_3_uop_decoded_branchCtrl_isIndirect;
    entries_3_uop_decoded_branchCtrl_laCfIdx <= entriesNext_3_uop_decoded_branchCtrl_laCfIdx;
    entries_3_uop_decoded_fpuCtrl_opType <= entriesNext_3_uop_decoded_fpuCtrl_opType;
    entries_3_uop_decoded_fpuCtrl_fpSizeSrc1 <= entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc1;
    entries_3_uop_decoded_fpuCtrl_fpSizeSrc2 <= entriesNext_3_uop_decoded_fpuCtrl_fpSizeSrc2;
    entries_3_uop_decoded_fpuCtrl_fpSizeDest <= entriesNext_3_uop_decoded_fpuCtrl_fpSizeDest;
    entries_3_uop_decoded_fpuCtrl_roundingMode <= entriesNext_3_uop_decoded_fpuCtrl_roundingMode;
    entries_3_uop_decoded_fpuCtrl_isIntegerDest <= entriesNext_3_uop_decoded_fpuCtrl_isIntegerDest;
    entries_3_uop_decoded_fpuCtrl_isSignedCvt <= entriesNext_3_uop_decoded_fpuCtrl_isSignedCvt;
    entries_3_uop_decoded_fpuCtrl_fmaNegSrc1 <= entriesNext_3_uop_decoded_fpuCtrl_fmaNegSrc1;
    entries_3_uop_decoded_fpuCtrl_fcmpCond <= entriesNext_3_uop_decoded_fpuCtrl_fcmpCond;
    entries_3_uop_decoded_csrCtrl_csrAddr <= entriesNext_3_uop_decoded_csrCtrl_csrAddr;
    entries_3_uop_decoded_csrCtrl_isWrite <= entriesNext_3_uop_decoded_csrCtrl_isWrite;
    entries_3_uop_decoded_csrCtrl_isRead <= entriesNext_3_uop_decoded_csrCtrl_isRead;
    entries_3_uop_decoded_csrCtrl_isExchange <= entriesNext_3_uop_decoded_csrCtrl_isExchange;
    entries_3_uop_decoded_csrCtrl_useUimmAsSrc <= entriesNext_3_uop_decoded_csrCtrl_useUimmAsSrc;
    entries_3_uop_decoded_sysCtrl_sysCode <= entriesNext_3_uop_decoded_sysCtrl_sysCode;
    entries_3_uop_decoded_sysCtrl_isExceptionReturn <= entriesNext_3_uop_decoded_sysCtrl_isExceptionReturn;
    entries_3_uop_decoded_sysCtrl_isTlbOp <= entriesNext_3_uop_decoded_sysCtrl_isTlbOp;
    entries_3_uop_decoded_sysCtrl_tlbOpType <= entriesNext_3_uop_decoded_sysCtrl_tlbOpType;
    entries_3_uop_decoded_decodeExceptionCode <= entriesNext_3_uop_decoded_decodeExceptionCode;
    entries_3_uop_decoded_hasDecodeException <= entriesNext_3_uop_decoded_hasDecodeException;
    entries_3_uop_decoded_isMicrocode <= entriesNext_3_uop_decoded_isMicrocode;
    entries_3_uop_decoded_microcodeEntry <= entriesNext_3_uop_decoded_microcodeEntry;
    entries_3_uop_decoded_isSerializing <= entriesNext_3_uop_decoded_isSerializing;
    entries_3_uop_decoded_isBranchOrJump <= entriesNext_3_uop_decoded_isBranchOrJump;
    entries_3_uop_decoded_branchPrediction_isTaken <= entriesNext_3_uop_decoded_branchPrediction_isTaken;
    entries_3_uop_decoded_branchPrediction_target <= entriesNext_3_uop_decoded_branchPrediction_target;
    entries_3_uop_decoded_branchPrediction_wasPredicted <= entriesNext_3_uop_decoded_branchPrediction_wasPredicted;
    entries_3_uop_rename_physSrc1_idx <= entriesNext_3_uop_rename_physSrc1_idx;
    entries_3_uop_rename_physSrc1IsFpr <= entriesNext_3_uop_rename_physSrc1IsFpr;
    entries_3_uop_rename_physSrc2_idx <= entriesNext_3_uop_rename_physSrc2_idx;
    entries_3_uop_rename_physSrc2IsFpr <= entriesNext_3_uop_rename_physSrc2IsFpr;
    entries_3_uop_rename_physDest_idx <= entriesNext_3_uop_rename_physDest_idx;
    entries_3_uop_rename_physDestIsFpr <= entriesNext_3_uop_rename_physDestIsFpr;
    entries_3_uop_rename_oldPhysDest_idx <= entriesNext_3_uop_rename_oldPhysDest_idx;
    entries_3_uop_rename_oldPhysDestIsFpr <= entriesNext_3_uop_rename_oldPhysDestIsFpr;
    entries_3_uop_rename_allocatesPhysDest <= entriesNext_3_uop_rename_allocatesPhysDest;
    entries_3_uop_rename_writesToPhysReg <= entriesNext_3_uop_rename_writesToPhysReg;
    entries_3_uop_robPtr <= entriesNext_3_uop_robPtr;
    entries_3_uop_uniqueId <= entriesNext_3_uop_uniqueId;
    entries_3_uop_dispatched <= entriesNext_3_uop_dispatched;
    entries_3_uop_executed <= entriesNext_3_uop_executed;
    entries_3_uop_hasException <= entriesNext_3_uop_hasException;
    entries_3_uop_exceptionCode <= entriesNext_3_uop_exceptionCode;
    entries_3_robPtr <= entriesNext_3_robPtr;
    entries_3_physDest_idx <= entriesNext_3_physDest_idx;
    entries_3_physDestIsFpr <= entriesNext_3_physDestIsFpr;
    entries_3_writesToPhysReg <= entriesNext_3_writesToPhysReg;
    entries_3_useSrc1 <= entriesNext_3_useSrc1;
    entries_3_src1Data <= entriesNext_3_src1Data;
    entries_3_src1Tag <= entriesNext_3_src1Tag;
    entries_3_src1Ready <= entriesNext_3_src1Ready;
    entries_3_src1IsFpr <= entriesNext_3_src1IsFpr;
    entries_3_useSrc2 <= entriesNext_3_useSrc2;
    entries_3_src2Data <= entriesNext_3_src2Data;
    entries_3_src2Tag <= entriesNext_3_src2Tag;
    entries_3_src2Ready <= entriesNext_3_src2Ready;
    entries_3_src2IsFpr <= entriesNext_3_src2IsFpr;
    entries_3_mulDivCtrl_valid <= entriesNext_3_mulDivCtrl_valid;
    entries_3_mulDivCtrl_isDiv <= entriesNext_3_mulDivCtrl_isDiv;
    entries_3_mulDivCtrl_isSigned <= entriesNext_3_mulDivCtrl_isSigned;
    entries_3_mulDivCtrl_isWordOp <= entriesNext_3_mulDivCtrl_isWordOp;
  end


endmodule

module IssueQueueComponent (
  input  wire          io_allocateIn_valid,
  output wire          io_allocateIn_ready,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_pc,
  input  wire          io_allocateIn_payload_uop_decoded_isValid,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_uopCode,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_exeUnit,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_isa,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archDest_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archDest_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_writeArchDestEn,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archSrc1_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archSrc1_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_useArchSrc1,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_archSrc2_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_archSrc2_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_useArchSrc2,
  input  wire          io_allocateIn_payload_uop_decoded_usePcForAddr,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_imm,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_immUsage,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isSub,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isAdd,
  input  wire          io_allocateIn_payload_uop_decoded_aluCtrl_isSigned,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_aluCtrl_logicOp,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isRight,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate,
  input  wire          io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_valid,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isDiv,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isSigned,
  input  wire          io_allocateIn_payload_uop_decoded_mulDivCtrl_isWordOp,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_memCtrl_size,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isSignedLoad,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isStore,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isLoadLinked,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isStoreCond,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_memCtrl_atomicOp,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isFence,
  input  wire [7:0]    io_allocateIn_payload_uop_decoded_memCtrl_fenceMode,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isCacheOp,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_memCtrl_cacheOpType,
  input  wire          io_allocateIn_payload_uop_decoded_memCtrl_isPrefetch,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_branchCtrl_condition,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isJump,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isLink,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_idx,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype,
  input  wire          io_allocateIn_payload_uop_decoded_branchCtrl_isIndirect,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_branchCtrl_laCfIdx,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_opType,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest,
  input  wire [2:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_roundingMode,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_isIntegerDest,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_isSignedCvt,
  input  wire          io_allocateIn_payload_uop_decoded_fpuCtrl_fmaNegSrc1,
  input  wire [4:0]    io_allocateIn_payload_uop_decoded_fpuCtrl_fcmpCond,
  input  wire [13:0]   io_allocateIn_payload_uop_decoded_csrCtrl_csrAddr,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isWrite,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isRead,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_isExchange,
  input  wire          io_allocateIn_payload_uop_decoded_csrCtrl_useUimmAsSrc,
  input  wire [19:0]   io_allocateIn_payload_uop_decoded_sysCtrl_sysCode,
  input  wire          io_allocateIn_payload_uop_decoded_sysCtrl_isExceptionReturn,
  input  wire          io_allocateIn_payload_uop_decoded_sysCtrl_isTlbOp,
  input  wire [3:0]    io_allocateIn_payload_uop_decoded_sysCtrl_tlbOpType,
  input  wire [1:0]    io_allocateIn_payload_uop_decoded_decodeExceptionCode,
  input  wire          io_allocateIn_payload_uop_decoded_hasDecodeException,
  input  wire          io_allocateIn_payload_uop_decoded_isMicrocode,
  input  wire [7:0]    io_allocateIn_payload_uop_decoded_microcodeEntry,
  input  wire          io_allocateIn_payload_uop_decoded_isSerializing,
  input  wire          io_allocateIn_payload_uop_decoded_isBranchOrJump,
  input  wire          io_allocateIn_payload_uop_decoded_branchPrediction_isTaken,
  input  wire [31:0]   io_allocateIn_payload_uop_decoded_branchPrediction_target,
  input  wire          io_allocateIn_payload_uop_decoded_branchPrediction_wasPredicted,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physSrc1_idx,
  input  wire          io_allocateIn_payload_uop_rename_physSrc1IsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physSrc2_idx,
  input  wire          io_allocateIn_payload_uop_rename_physSrc2IsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_physDest_idx,
  input  wire          io_allocateIn_payload_uop_rename_physDestIsFpr,
  input  wire [5:0]    io_allocateIn_payload_uop_rename_oldPhysDest_idx,
  input  wire          io_allocateIn_payload_uop_rename_oldPhysDestIsFpr,
  input  wire          io_allocateIn_payload_uop_rename_allocatesPhysDest,
  input  wire          io_allocateIn_payload_uop_rename_writesToPhysReg,
  input  wire [3:0]    io_allocateIn_payload_uop_robPtr,
  input  wire [15:0]   io_allocateIn_payload_uop_uniqueId,
  input  wire          io_allocateIn_payload_uop_dispatched,
  input  wire          io_allocateIn_payload_uop_executed,
  input  wire          io_allocateIn_payload_uop_hasException,
  input  wire [7:0]    io_allocateIn_payload_uop_exceptionCode,
  input  wire          io_allocateIn_payload_src1InitialReady,
  input  wire          io_allocateIn_payload_src2InitialReady,
  output wire          io_issueOut_valid,
  input  wire          io_issueOut_ready,
  output wire [3:0]    io_issueOut_payload_robPtr,
  output wire [5:0]    io_issueOut_payload_physDest_idx,
  output wire          io_issueOut_payload_physDestIsFpr,
  output wire          io_issueOut_payload_writesToPhysReg,
  output wire          io_issueOut_payload_useSrc1,
  output wire [31:0]   io_issueOut_payload_src1Data,
  output wire [5:0]    io_issueOut_payload_src1Tag,
  output wire          io_issueOut_payload_src1Ready,
  output wire          io_issueOut_payload_src1IsFpr,
  output wire          io_issueOut_payload_useSrc2,
  output wire [31:0]   io_issueOut_payload_src2Data,
  output wire [5:0]    io_issueOut_payload_src2Tag,
  output wire          io_issueOut_payload_src2Ready,
  output wire          io_issueOut_payload_src2IsFpr,
  output wire          io_issueOut_payload_aluCtrl_valid,
  output wire          io_issueOut_payload_aluCtrl_isSub,
  output wire          io_issueOut_payload_aluCtrl_isAdd,
  output wire          io_issueOut_payload_aluCtrl_isSigned,
  output wire [1:0]    io_issueOut_payload_aluCtrl_logicOp,
  output wire          io_issueOut_payload_shiftCtrl_valid,
  output wire          io_issueOut_payload_shiftCtrl_isRight,
  output wire          io_issueOut_payload_shiftCtrl_isArithmetic,
  output wire          io_issueOut_payload_shiftCtrl_isRotate,
  output wire          io_issueOut_payload_shiftCtrl_isDoubleWord,
  output wire [31:0]   io_issueOut_payload_imm,
  output wire [2:0]    io_issueOut_payload_immUsage,
  input  wire          io_wakeupIn_0_valid,
  input  wire [5:0]    io_wakeupIn_0_payload_physRegIdx,
  input  wire          io_wakeupIn_1_valid,
  input  wire [5:0]    io_wakeupIn_1_payload_physRegIdx,
  input  wire          io_wakeupIn_2_valid,
  input  wire [5:0]    io_wakeupIn_2_payload_physRegIdx,
  input  wire          io_wakeupIn_3_valid,
  input  wire [5:0]    io_wakeupIn_3_payload_physRegIdx,
  input  wire          io_wakeupIn_4_valid,
  input  wire [5:0]    io_wakeupIn_4_payload_physRegIdx,
  input  wire          io_flush,
  input  wire          clk,
  input  wire          reset
);
  localparam BaseUopCode_NOP = 5'd0;
  localparam BaseUopCode_ILLEGAL = 5'd1;
  localparam BaseUopCode_ALU = 5'd2;
  localparam BaseUopCode_SHIFT = 5'd3;
  localparam BaseUopCode_MUL = 5'd4;
  localparam BaseUopCode_DIV = 5'd5;
  localparam BaseUopCode_LOAD = 5'd6;
  localparam BaseUopCode_STORE = 5'd7;
  localparam BaseUopCode_ATOMIC = 5'd8;
  localparam BaseUopCode_MEM_BARRIER = 5'd9;
  localparam BaseUopCode_PREFETCH = 5'd10;
  localparam BaseUopCode_BRANCH = 5'd11;
  localparam BaseUopCode_JUMP_REG = 5'd12;
  localparam BaseUopCode_JUMP_IMM = 5'd13;
  localparam BaseUopCode_SYSTEM_OP = 5'd14;
  localparam BaseUopCode_CSR_ACCESS = 5'd15;
  localparam BaseUopCode_FPU_ALU = 5'd16;
  localparam BaseUopCode_FPU_CVT = 5'd17;
  localparam BaseUopCode_FPU_CMP = 5'd18;
  localparam BaseUopCode_FPU_SEL = 5'd19;
  localparam BaseUopCode_LA_BITMANIP = 5'd20;
  localparam BaseUopCode_LA_CACOP = 5'd21;
  localparam BaseUopCode_LA_TLB = 5'd22;
  localparam BaseUopCode_IDLE = 5'd23;
  localparam ExeUnitType_NONE = 4'd0;
  localparam ExeUnitType_ALU_INT = 4'd1;
  localparam ExeUnitType_MUL_INT = 4'd2;
  localparam ExeUnitType_DIV_INT = 4'd3;
  localparam ExeUnitType_MEM = 4'd4;
  localparam ExeUnitType_BRU = 4'd5;
  localparam ExeUnitType_CSR = 4'd6;
  localparam ExeUnitType_FPU_ADD_MUL_CVT_CMP = 4'd7;
  localparam ExeUnitType_FPU_DIV_SQRT = 4'd8;
  localparam IsaType_UNKNOWN = 2'd0;
  localparam IsaType_DEMO = 2'd1;
  localparam IsaType_RISCV = 2'd2;
  localparam IsaType_LOONGARCH = 2'd3;
  localparam ArchRegType_GPR = 2'd0;
  localparam ArchRegType_FPR = 2'd1;
  localparam ArchRegType_CSR = 2'd2;
  localparam ArchRegType_LA_CF = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;
  localparam BranchCondition_NUL = 5'd0;
  localparam BranchCondition_EQ = 5'd1;
  localparam BranchCondition_NE = 5'd2;
  localparam BranchCondition_LT = 5'd3;
  localparam BranchCondition_GE = 5'd4;
  localparam BranchCondition_LTU = 5'd5;
  localparam BranchCondition_GEU = 5'd6;
  localparam BranchCondition_EQZ = 5'd7;
  localparam BranchCondition_NEZ = 5'd8;
  localparam BranchCondition_LTZ = 5'd9;
  localparam BranchCondition_GEZ = 5'd10;
  localparam BranchCondition_GTZ = 5'd11;
  localparam BranchCondition_LEZ = 5'd12;
  localparam BranchCondition_F_EQ = 5'd13;
  localparam BranchCondition_F_NE = 5'd14;
  localparam BranchCondition_F_LT = 5'd15;
  localparam BranchCondition_F_LE = 5'd16;
  localparam BranchCondition_F_UN = 5'd17;
  localparam BranchCondition_LA_CF_TRUE = 5'd18;
  localparam BranchCondition_LA_CF_FALSE = 5'd19;
  localparam DecodeExCode_INVALID = 2'd0;
  localparam DecodeExCode_FETCH_ERROR = 2'd1;
  localparam DecodeExCode_DECODE_ERROR = 2'd2;
  localparam DecodeExCode_OK = 2'd3;

  wire       [3:0]    _zz_issueRequestMask_ohFirst_masked;
  reg        [1:0]    _zz__zz_io_issueOut_payload_aluCtrl_logicOp;
  reg        [2:0]    _zz__zz_io_issueOut_payload_immUsage;
  reg        [3:0]    _zz_io_issueOut_payload_robPtr;
  reg        [5:0]    _zz_io_issueOut_payload_physDest_idx;
  reg                 _zz_io_issueOut_payload_physDestIsFpr;
  reg                 _zz_io_issueOut_payload_writesToPhysReg;
  reg                 _zz_io_issueOut_payload_useSrc1;
  reg        [31:0]   _zz_io_issueOut_payload_src1Data;
  reg        [5:0]    _zz_io_issueOut_payload_src1Tag;
  reg                 _zz_io_issueOut_payload_src1Ready;
  reg                 _zz_io_issueOut_payload_src1IsFpr;
  reg                 _zz_io_issueOut_payload_useSrc2;
  reg        [31:0]   _zz_io_issueOut_payload_src2Data;
  reg        [5:0]    _zz_io_issueOut_payload_src2Tag;
  reg                 _zz_io_issueOut_payload_src2Ready;
  reg                 _zz_io_issueOut_payload_src2IsFpr;
  reg                 _zz_io_issueOut_payload_aluCtrl_valid;
  reg                 _zz_io_issueOut_payload_aluCtrl_isSub;
  reg                 _zz_io_issueOut_payload_aluCtrl_isAdd;
  reg                 _zz_io_issueOut_payload_aluCtrl_isSigned;
  reg                 _zz_io_issueOut_payload_shiftCtrl_valid;
  reg                 _zz_io_issueOut_payload_shiftCtrl_isRight;
  reg                 _zz_io_issueOut_payload_shiftCtrl_isArithmetic;
  reg                 _zz_io_issueOut_payload_shiftCtrl_isRotate;
  reg                 _zz_io_issueOut_payload_shiftCtrl_isDoubleWord;
  reg        [31:0]   _zz_io_issueOut_payload_imm;
  wire       [3:0]    _zz_allocationMask_1;
  reg        [2:0]    _zz_currentValidCount_8;
  wire       [2:0]    _zz_currentValidCount_9;
  reg        [2:0]    _zz_currentValidCount_10;
  wire       [2:0]    _zz_currentValidCount_11;
  wire       [0:0]    _zz_currentValidCount_12;
  reg        [3:0]    entries_0_robPtr;
  reg        [5:0]    entries_0_physDest_idx;
  reg                 entries_0_physDestIsFpr;
  reg                 entries_0_writesToPhysReg;
  reg                 entries_0_useSrc1;
  reg        [31:0]   entries_0_src1Data;
  reg        [5:0]    entries_0_src1Tag;
  reg                 entries_0_src1Ready;
  reg                 entries_0_src1IsFpr;
  reg                 entries_0_useSrc2;
  reg        [31:0]   entries_0_src2Data;
  reg        [5:0]    entries_0_src2Tag;
  reg                 entries_0_src2Ready;
  reg                 entries_0_src2IsFpr;
  reg                 entries_0_aluCtrl_valid;
  reg                 entries_0_aluCtrl_isSub;
  reg                 entries_0_aluCtrl_isAdd;
  reg                 entries_0_aluCtrl_isSigned;
  reg        [1:0]    entries_0_aluCtrl_logicOp;
  reg                 entries_0_shiftCtrl_valid;
  reg                 entries_0_shiftCtrl_isRight;
  reg                 entries_0_shiftCtrl_isArithmetic;
  reg                 entries_0_shiftCtrl_isRotate;
  reg                 entries_0_shiftCtrl_isDoubleWord;
  reg        [31:0]   entries_0_imm;
  reg        [2:0]    entries_0_immUsage;
  reg        [3:0]    entries_1_robPtr;
  reg        [5:0]    entries_1_physDest_idx;
  reg                 entries_1_physDestIsFpr;
  reg                 entries_1_writesToPhysReg;
  reg                 entries_1_useSrc1;
  reg        [31:0]   entries_1_src1Data;
  reg        [5:0]    entries_1_src1Tag;
  reg                 entries_1_src1Ready;
  reg                 entries_1_src1IsFpr;
  reg                 entries_1_useSrc2;
  reg        [31:0]   entries_1_src2Data;
  reg        [5:0]    entries_1_src2Tag;
  reg                 entries_1_src2Ready;
  reg                 entries_1_src2IsFpr;
  reg                 entries_1_aluCtrl_valid;
  reg                 entries_1_aluCtrl_isSub;
  reg                 entries_1_aluCtrl_isAdd;
  reg                 entries_1_aluCtrl_isSigned;
  reg        [1:0]    entries_1_aluCtrl_logicOp;
  reg                 entries_1_shiftCtrl_valid;
  reg                 entries_1_shiftCtrl_isRight;
  reg                 entries_1_shiftCtrl_isArithmetic;
  reg                 entries_1_shiftCtrl_isRotate;
  reg                 entries_1_shiftCtrl_isDoubleWord;
  reg        [31:0]   entries_1_imm;
  reg        [2:0]    entries_1_immUsage;
  reg        [3:0]    entries_2_robPtr;
  reg        [5:0]    entries_2_physDest_idx;
  reg                 entries_2_physDestIsFpr;
  reg                 entries_2_writesToPhysReg;
  reg                 entries_2_useSrc1;
  reg        [31:0]   entries_2_src1Data;
  reg        [5:0]    entries_2_src1Tag;
  reg                 entries_2_src1Ready;
  reg                 entries_2_src1IsFpr;
  reg                 entries_2_useSrc2;
  reg        [31:0]   entries_2_src2Data;
  reg        [5:0]    entries_2_src2Tag;
  reg                 entries_2_src2Ready;
  reg                 entries_2_src2IsFpr;
  reg                 entries_2_aluCtrl_valid;
  reg                 entries_2_aluCtrl_isSub;
  reg                 entries_2_aluCtrl_isAdd;
  reg                 entries_2_aluCtrl_isSigned;
  reg        [1:0]    entries_2_aluCtrl_logicOp;
  reg                 entries_2_shiftCtrl_valid;
  reg                 entries_2_shiftCtrl_isRight;
  reg                 entries_2_shiftCtrl_isArithmetic;
  reg                 entries_2_shiftCtrl_isRotate;
  reg                 entries_2_shiftCtrl_isDoubleWord;
  reg        [31:0]   entries_2_imm;
  reg        [2:0]    entries_2_immUsage;
  reg        [3:0]    entries_3_robPtr;
  reg        [5:0]    entries_3_physDest_idx;
  reg                 entries_3_physDestIsFpr;
  reg                 entries_3_writesToPhysReg;
  reg                 entries_3_useSrc1;
  reg        [31:0]   entries_3_src1Data;
  reg        [5:0]    entries_3_src1Tag;
  reg                 entries_3_src1Ready;
  reg                 entries_3_src1IsFpr;
  reg                 entries_3_useSrc2;
  reg        [31:0]   entries_3_src2Data;
  reg        [5:0]    entries_3_src2Tag;
  reg                 entries_3_src2Ready;
  reg                 entries_3_src2IsFpr;
  reg                 entries_3_aluCtrl_valid;
  reg                 entries_3_aluCtrl_isSub;
  reg                 entries_3_aluCtrl_isAdd;
  reg                 entries_3_aluCtrl_isSigned;
  reg        [1:0]    entries_3_aluCtrl_logicOp;
  reg                 entries_3_shiftCtrl_valid;
  reg                 entries_3_shiftCtrl_isRight;
  reg                 entries_3_shiftCtrl_isArithmetic;
  reg                 entries_3_shiftCtrl_isRotate;
  reg                 entries_3_shiftCtrl_isDoubleWord;
  reg        [31:0]   entries_3_imm;
  reg        [2:0]    entries_3_immUsage;
  reg                 entryValids_0;
  reg                 entryValids_1;
  reg                 entryValids_2;
  reg                 entryValids_3;
  wire                io_issueOut_fire;
  wire                localWakeupValid;
  reg        [3:0]    wokeUpSrc1Mask;
  reg        [3:0]    wokeUpSrc2Mask;
  wire                _zz_when_IssueQueueComponent_l103;
  wire                _zz_when_IssueQueueComponent_l106;
  wire                when_IssueQueueComponent_l103;
  wire                when_IssueQueueComponent_l106;
  wire                when_IssueQueueComponent_l113;
  wire                when_IssueQueueComponent_l116;
  wire                when_IssueQueueComponent_l113_1;
  wire                when_IssueQueueComponent_l116_1;
  wire                when_IssueQueueComponent_l113_2;
  wire                when_IssueQueueComponent_l116_2;
  wire                when_IssueQueueComponent_l113_3;
  wire                when_IssueQueueComponent_l116_3;
  wire                when_IssueQueueComponent_l113_4;
  wire                when_IssueQueueComponent_l116_4;
  wire                _zz_when_IssueQueueComponent_l103_1;
  wire                _zz_when_IssueQueueComponent_l106_1;
  wire                when_IssueQueueComponent_l103_1;
  wire                when_IssueQueueComponent_l106_1;
  wire                when_IssueQueueComponent_l113_5;
  wire                when_IssueQueueComponent_l116_5;
  wire                when_IssueQueueComponent_l113_6;
  wire                when_IssueQueueComponent_l116_6;
  wire                when_IssueQueueComponent_l113_7;
  wire                when_IssueQueueComponent_l116_7;
  wire                when_IssueQueueComponent_l113_8;
  wire                when_IssueQueueComponent_l116_8;
  wire                when_IssueQueueComponent_l113_9;
  wire                when_IssueQueueComponent_l116_9;
  wire                _zz_when_IssueQueueComponent_l103_2;
  wire                _zz_when_IssueQueueComponent_l106_2;
  wire                when_IssueQueueComponent_l103_2;
  wire                when_IssueQueueComponent_l106_2;
  wire                when_IssueQueueComponent_l113_10;
  wire                when_IssueQueueComponent_l116_10;
  wire                when_IssueQueueComponent_l113_11;
  wire                when_IssueQueueComponent_l116_11;
  wire                when_IssueQueueComponent_l113_12;
  wire                when_IssueQueueComponent_l116_12;
  wire                when_IssueQueueComponent_l113_13;
  wire                when_IssueQueueComponent_l116_13;
  wire                when_IssueQueueComponent_l113_14;
  wire                when_IssueQueueComponent_l116_14;
  wire                _zz_when_IssueQueueComponent_l103_3;
  wire                _zz_when_IssueQueueComponent_l106_3;
  wire                when_IssueQueueComponent_l103_3;
  wire                when_IssueQueueComponent_l106_3;
  wire                when_IssueQueueComponent_l113_15;
  wire                when_IssueQueueComponent_l116_15;
  wire                when_IssueQueueComponent_l113_16;
  wire                when_IssueQueueComponent_l116_16;
  wire                when_IssueQueueComponent_l113_17;
  wire                when_IssueQueueComponent_l116_17;
  wire                when_IssueQueueComponent_l113_18;
  wire                when_IssueQueueComponent_l116_18;
  wire                when_IssueQueueComponent_l113_19;
  wire                when_IssueQueueComponent_l116_19;
  wire                entriesReadyToIssue_0;
  wire                entriesReadyToIssue_1;
  wire                entriesReadyToIssue_2;
  wire                entriesReadyToIssue_3;
  wire       [3:0]    issueRequestMask;
  wire       [3:0]    issueRequestMask_ohFirst_input;
  wire       [3:0]    issueRequestMask_ohFirst_masked;
  wire       [3:0]    issueRequestOh;
  wire                _zz_issueIdx;
  wire                _zz_issueIdx_1;
  wire                _zz_issueIdx_2;
  wire       [1:0]    issueIdx;
  wire       [1:0]    _zz_io_issueOut_payload_aluCtrl_logicOp;
  wire       [2:0]    _zz_io_issueOut_payload_immUsage;
  wire       [3:0]    freeSlotsMask;
  wire                hasSpaceForNewEntry;
  reg        [3:0]    firedSlotMask;
  wire       [3:0]    _zz_allocationMask;
  wire       [3:0]    allocationMask;
  wire                _zz_allocateIdx;
  wire                _zz_allocateIdx_1;
  wire                _zz_allocateIdx_2;
  wire       [1:0]    allocateIdx;
  reg        [3:0]    entriesNext_0_robPtr;
  reg        [5:0]    entriesNext_0_physDest_idx;
  reg                 entriesNext_0_physDestIsFpr;
  reg                 entriesNext_0_writesToPhysReg;
  reg                 entriesNext_0_useSrc1;
  reg        [31:0]   entriesNext_0_src1Data;
  reg        [5:0]    entriesNext_0_src1Tag;
  reg                 entriesNext_0_src1Ready;
  reg                 entriesNext_0_src1IsFpr;
  reg                 entriesNext_0_useSrc2;
  reg        [31:0]   entriesNext_0_src2Data;
  reg        [5:0]    entriesNext_0_src2Tag;
  reg                 entriesNext_0_src2Ready;
  reg                 entriesNext_0_src2IsFpr;
  reg                 entriesNext_0_aluCtrl_valid;
  reg                 entriesNext_0_aluCtrl_isSub;
  reg                 entriesNext_0_aluCtrl_isAdd;
  reg                 entriesNext_0_aluCtrl_isSigned;
  reg        [1:0]    entriesNext_0_aluCtrl_logicOp;
  reg                 entriesNext_0_shiftCtrl_valid;
  reg                 entriesNext_0_shiftCtrl_isRight;
  reg                 entriesNext_0_shiftCtrl_isArithmetic;
  reg                 entriesNext_0_shiftCtrl_isRotate;
  reg                 entriesNext_0_shiftCtrl_isDoubleWord;
  reg        [31:0]   entriesNext_0_imm;
  reg        [2:0]    entriesNext_0_immUsage;
  reg        [3:0]    entriesNext_1_robPtr;
  reg        [5:0]    entriesNext_1_physDest_idx;
  reg                 entriesNext_1_physDestIsFpr;
  reg                 entriesNext_1_writesToPhysReg;
  reg                 entriesNext_1_useSrc1;
  reg        [31:0]   entriesNext_1_src1Data;
  reg        [5:0]    entriesNext_1_src1Tag;
  reg                 entriesNext_1_src1Ready;
  reg                 entriesNext_1_src1IsFpr;
  reg                 entriesNext_1_useSrc2;
  reg        [31:0]   entriesNext_1_src2Data;
  reg        [5:0]    entriesNext_1_src2Tag;
  reg                 entriesNext_1_src2Ready;
  reg                 entriesNext_1_src2IsFpr;
  reg                 entriesNext_1_aluCtrl_valid;
  reg                 entriesNext_1_aluCtrl_isSub;
  reg                 entriesNext_1_aluCtrl_isAdd;
  reg                 entriesNext_1_aluCtrl_isSigned;
  reg        [1:0]    entriesNext_1_aluCtrl_logicOp;
  reg                 entriesNext_1_shiftCtrl_valid;
  reg                 entriesNext_1_shiftCtrl_isRight;
  reg                 entriesNext_1_shiftCtrl_isArithmetic;
  reg                 entriesNext_1_shiftCtrl_isRotate;
  reg                 entriesNext_1_shiftCtrl_isDoubleWord;
  reg        [31:0]   entriesNext_1_imm;
  reg        [2:0]    entriesNext_1_immUsage;
  reg        [3:0]    entriesNext_2_robPtr;
  reg        [5:0]    entriesNext_2_physDest_idx;
  reg                 entriesNext_2_physDestIsFpr;
  reg                 entriesNext_2_writesToPhysReg;
  reg                 entriesNext_2_useSrc1;
  reg        [31:0]   entriesNext_2_src1Data;
  reg        [5:0]    entriesNext_2_src1Tag;
  reg                 entriesNext_2_src1Ready;
  reg                 entriesNext_2_src1IsFpr;
  reg                 entriesNext_2_useSrc2;
  reg        [31:0]   entriesNext_2_src2Data;
  reg        [5:0]    entriesNext_2_src2Tag;
  reg                 entriesNext_2_src2Ready;
  reg                 entriesNext_2_src2IsFpr;
  reg                 entriesNext_2_aluCtrl_valid;
  reg                 entriesNext_2_aluCtrl_isSub;
  reg                 entriesNext_2_aluCtrl_isAdd;
  reg                 entriesNext_2_aluCtrl_isSigned;
  reg        [1:0]    entriesNext_2_aluCtrl_logicOp;
  reg                 entriesNext_2_shiftCtrl_valid;
  reg                 entriesNext_2_shiftCtrl_isRight;
  reg                 entriesNext_2_shiftCtrl_isArithmetic;
  reg                 entriesNext_2_shiftCtrl_isRotate;
  reg                 entriesNext_2_shiftCtrl_isDoubleWord;
  reg        [31:0]   entriesNext_2_imm;
  reg        [2:0]    entriesNext_2_immUsage;
  reg        [3:0]    entriesNext_3_robPtr;
  reg        [5:0]    entriesNext_3_physDest_idx;
  reg                 entriesNext_3_physDestIsFpr;
  reg                 entriesNext_3_writesToPhysReg;
  reg                 entriesNext_3_useSrc1;
  reg        [31:0]   entriesNext_3_src1Data;
  reg        [5:0]    entriesNext_3_src1Tag;
  reg                 entriesNext_3_src1Ready;
  reg                 entriesNext_3_src1IsFpr;
  reg                 entriesNext_3_useSrc2;
  reg        [31:0]   entriesNext_3_src2Data;
  reg        [5:0]    entriesNext_3_src2Tag;
  reg                 entriesNext_3_src2Ready;
  reg                 entriesNext_3_src2IsFpr;
  reg                 entriesNext_3_aluCtrl_valid;
  reg                 entriesNext_3_aluCtrl_isSub;
  reg                 entriesNext_3_aluCtrl_isAdd;
  reg                 entriesNext_3_aluCtrl_isSigned;
  reg        [1:0]    entriesNext_3_aluCtrl_logicOp;
  reg                 entriesNext_3_shiftCtrl_valid;
  reg                 entriesNext_3_shiftCtrl_isRight;
  reg                 entriesNext_3_shiftCtrl_isArithmetic;
  reg                 entriesNext_3_shiftCtrl_isRotate;
  reg                 entriesNext_3_shiftCtrl_isDoubleWord;
  reg        [31:0]   entriesNext_3_imm;
  reg        [2:0]    entriesNext_3_immUsage;
  reg                 entryValidsNext_0;
  reg                 entryValidsNext_1;
  reg                 entryValidsNext_2;
  reg                 entryValidsNext_3;
  wire                when_IssueQueueComponent_l186;
  wire                when_IssueQueueComponent_l187;
  wire                when_IssueQueueComponent_l186_1;
  wire                when_IssueQueueComponent_l187_1;
  wire                when_IssueQueueComponent_l186_2;
  wire                when_IssueQueueComponent_l187_2;
  wire                when_IssueQueueComponent_l186_3;
  wire                when_IssueQueueComponent_l187_3;
  wire       [3:0]    _zz_1;
  wire                io_allocateIn_fire;
  wire       [3:0]    _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_entriesNext_0_src1Ready;
  wire                _zz_entriesNext_0_src2Ready;
  wire       [3:0]    _zz_7;
  wire                when_IssueQueueComponent_l212;
  wire                when_IssueQueueComponent_l215;
  wire                when_IssueQueueComponent_l212_1;
  wire                when_IssueQueueComponent_l215_1;
  wire                when_IssueQueueComponent_l212_2;
  wire                when_IssueQueueComponent_l215_2;
  wire                when_IssueQueueComponent_l212_3;
  wire                when_IssueQueueComponent_l215_3;
  wire                when_IssueQueueComponent_l212_4;
  wire                when_IssueQueueComponent_l215_4;
  wire       [2:0]    _zz_currentValidCount;
  wire       [2:0]    _zz_currentValidCount_1;
  wire       [2:0]    _zz_currentValidCount_2;
  wire       [2:0]    _zz_currentValidCount_3;
  wire       [2:0]    _zz_currentValidCount_4;
  wire       [2:0]    _zz_currentValidCount_5;
  wire       [2:0]    _zz_currentValidCount_6;
  wire       [2:0]    _zz_currentValidCount_7;
  wire       [2:0]    currentValidCount;
  wire                logCondition;
  wire                when_IssueQueueComponent_l256;
  `ifndef SYNTHESIS
  reg [87:0] io_allocateIn_payload_uop_decoded_uopCode_string;
  reg [151:0] io_allocateIn_payload_uop_decoded_exeUnit_string;
  reg [71:0] io_allocateIn_payload_uop_decoded_isa_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] io_allocateIn_payload_uop_decoded_immUsage_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] io_allocateIn_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_allocateIn_payload_uop_decoded_decodeExceptionCode_string;
  reg [39:0] io_issueOut_payload_aluCtrl_logicOp_string;
  reg [103:0] io_issueOut_payload_immUsage_string;
  reg [39:0] entries_0_aluCtrl_logicOp_string;
  reg [103:0] entries_0_immUsage_string;
  reg [39:0] entries_1_aluCtrl_logicOp_string;
  reg [103:0] entries_1_immUsage_string;
  reg [39:0] entries_2_aluCtrl_logicOp_string;
  reg [103:0] entries_2_immUsage_string;
  reg [39:0] entries_3_aluCtrl_logicOp_string;
  reg [103:0] entries_3_immUsage_string;
  reg [39:0] _zz_io_issueOut_payload_aluCtrl_logicOp_string;
  reg [103:0] _zz_io_issueOut_payload_immUsage_string;
  reg [39:0] entriesNext_0_aluCtrl_logicOp_string;
  reg [103:0] entriesNext_0_immUsage_string;
  reg [39:0] entriesNext_1_aluCtrl_logicOp_string;
  reg [103:0] entriesNext_1_immUsage_string;
  reg [39:0] entriesNext_2_aluCtrl_logicOp_string;
  reg [103:0] entriesNext_2_immUsage_string;
  reg [39:0] entriesNext_3_aluCtrl_logicOp_string;
  reg [103:0] entriesNext_3_immUsage_string;
  `endif


  assign _zz_issueRequestMask_ohFirst_masked = (issueRequestMask_ohFirst_input - 4'b0001);
  assign _zz_allocationMask_1 = (_zz_allocationMask - 4'b0001);
  assign _zz_currentValidCount_12 = entryValids_3;
  assign _zz_currentValidCount_11 = {2'd0, _zz_currentValidCount_12};
  assign _zz_currentValidCount_9 = {entryValids_2,{entryValids_1,entryValids_0}};
  always @(*) begin
    case(issueIdx)
      2'b00 : begin
        _zz__zz_io_issueOut_payload_aluCtrl_logicOp = entries_0_aluCtrl_logicOp;
        _zz__zz_io_issueOut_payload_immUsage = entries_0_immUsage;
        _zz_io_issueOut_payload_robPtr = entries_0_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_0_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_0_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_0_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_0_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_0_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_0_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_0_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_0_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_0_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_0_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_0_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_0_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_0_src2IsFpr;
        _zz_io_issueOut_payload_aluCtrl_valid = entries_0_aluCtrl_valid;
        _zz_io_issueOut_payload_aluCtrl_isSub = entries_0_aluCtrl_isSub;
        _zz_io_issueOut_payload_aluCtrl_isAdd = entries_0_aluCtrl_isAdd;
        _zz_io_issueOut_payload_aluCtrl_isSigned = entries_0_aluCtrl_isSigned;
        _zz_io_issueOut_payload_shiftCtrl_valid = entries_0_shiftCtrl_valid;
        _zz_io_issueOut_payload_shiftCtrl_isRight = entries_0_shiftCtrl_isRight;
        _zz_io_issueOut_payload_shiftCtrl_isArithmetic = entries_0_shiftCtrl_isArithmetic;
        _zz_io_issueOut_payload_shiftCtrl_isRotate = entries_0_shiftCtrl_isRotate;
        _zz_io_issueOut_payload_shiftCtrl_isDoubleWord = entries_0_shiftCtrl_isDoubleWord;
        _zz_io_issueOut_payload_imm = entries_0_imm;
      end
      2'b01 : begin
        _zz__zz_io_issueOut_payload_aluCtrl_logicOp = entries_1_aluCtrl_logicOp;
        _zz__zz_io_issueOut_payload_immUsage = entries_1_immUsage;
        _zz_io_issueOut_payload_robPtr = entries_1_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_1_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_1_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_1_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_1_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_1_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_1_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_1_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_1_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_1_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_1_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_1_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_1_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_1_src2IsFpr;
        _zz_io_issueOut_payload_aluCtrl_valid = entries_1_aluCtrl_valid;
        _zz_io_issueOut_payload_aluCtrl_isSub = entries_1_aluCtrl_isSub;
        _zz_io_issueOut_payload_aluCtrl_isAdd = entries_1_aluCtrl_isAdd;
        _zz_io_issueOut_payload_aluCtrl_isSigned = entries_1_aluCtrl_isSigned;
        _zz_io_issueOut_payload_shiftCtrl_valid = entries_1_shiftCtrl_valid;
        _zz_io_issueOut_payload_shiftCtrl_isRight = entries_1_shiftCtrl_isRight;
        _zz_io_issueOut_payload_shiftCtrl_isArithmetic = entries_1_shiftCtrl_isArithmetic;
        _zz_io_issueOut_payload_shiftCtrl_isRotate = entries_1_shiftCtrl_isRotate;
        _zz_io_issueOut_payload_shiftCtrl_isDoubleWord = entries_1_shiftCtrl_isDoubleWord;
        _zz_io_issueOut_payload_imm = entries_1_imm;
      end
      2'b10 : begin
        _zz__zz_io_issueOut_payload_aluCtrl_logicOp = entries_2_aluCtrl_logicOp;
        _zz__zz_io_issueOut_payload_immUsage = entries_2_immUsage;
        _zz_io_issueOut_payload_robPtr = entries_2_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_2_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_2_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_2_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_2_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_2_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_2_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_2_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_2_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_2_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_2_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_2_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_2_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_2_src2IsFpr;
        _zz_io_issueOut_payload_aluCtrl_valid = entries_2_aluCtrl_valid;
        _zz_io_issueOut_payload_aluCtrl_isSub = entries_2_aluCtrl_isSub;
        _zz_io_issueOut_payload_aluCtrl_isAdd = entries_2_aluCtrl_isAdd;
        _zz_io_issueOut_payload_aluCtrl_isSigned = entries_2_aluCtrl_isSigned;
        _zz_io_issueOut_payload_shiftCtrl_valid = entries_2_shiftCtrl_valid;
        _zz_io_issueOut_payload_shiftCtrl_isRight = entries_2_shiftCtrl_isRight;
        _zz_io_issueOut_payload_shiftCtrl_isArithmetic = entries_2_shiftCtrl_isArithmetic;
        _zz_io_issueOut_payload_shiftCtrl_isRotate = entries_2_shiftCtrl_isRotate;
        _zz_io_issueOut_payload_shiftCtrl_isDoubleWord = entries_2_shiftCtrl_isDoubleWord;
        _zz_io_issueOut_payload_imm = entries_2_imm;
      end
      default : begin
        _zz__zz_io_issueOut_payload_aluCtrl_logicOp = entries_3_aluCtrl_logicOp;
        _zz__zz_io_issueOut_payload_immUsage = entries_3_immUsage;
        _zz_io_issueOut_payload_robPtr = entries_3_robPtr;
        _zz_io_issueOut_payload_physDest_idx = entries_3_physDest_idx;
        _zz_io_issueOut_payload_physDestIsFpr = entries_3_physDestIsFpr;
        _zz_io_issueOut_payload_writesToPhysReg = entries_3_writesToPhysReg;
        _zz_io_issueOut_payload_useSrc1 = entries_3_useSrc1;
        _zz_io_issueOut_payload_src1Data = entries_3_src1Data;
        _zz_io_issueOut_payload_src1Tag = entries_3_src1Tag;
        _zz_io_issueOut_payload_src1Ready = entries_3_src1Ready;
        _zz_io_issueOut_payload_src1IsFpr = entries_3_src1IsFpr;
        _zz_io_issueOut_payload_useSrc2 = entries_3_useSrc2;
        _zz_io_issueOut_payload_src2Data = entries_3_src2Data;
        _zz_io_issueOut_payload_src2Tag = entries_3_src2Tag;
        _zz_io_issueOut_payload_src2Ready = entries_3_src2Ready;
        _zz_io_issueOut_payload_src2IsFpr = entries_3_src2IsFpr;
        _zz_io_issueOut_payload_aluCtrl_valid = entries_3_aluCtrl_valid;
        _zz_io_issueOut_payload_aluCtrl_isSub = entries_3_aluCtrl_isSub;
        _zz_io_issueOut_payload_aluCtrl_isAdd = entries_3_aluCtrl_isAdd;
        _zz_io_issueOut_payload_aluCtrl_isSigned = entries_3_aluCtrl_isSigned;
        _zz_io_issueOut_payload_shiftCtrl_valid = entries_3_shiftCtrl_valid;
        _zz_io_issueOut_payload_shiftCtrl_isRight = entries_3_shiftCtrl_isRight;
        _zz_io_issueOut_payload_shiftCtrl_isArithmetic = entries_3_shiftCtrl_isArithmetic;
        _zz_io_issueOut_payload_shiftCtrl_isRotate = entries_3_shiftCtrl_isRotate;
        _zz_io_issueOut_payload_shiftCtrl_isDoubleWord = entries_3_shiftCtrl_isDoubleWord;
        _zz_io_issueOut_payload_imm = entries_3_imm;
      end
    endcase
  end

  always @(*) begin
    case(_zz_currentValidCount_9)
      3'b000 : _zz_currentValidCount_8 = _zz_currentValidCount;
      3'b001 : _zz_currentValidCount_8 = _zz_currentValidCount_1;
      3'b010 : _zz_currentValidCount_8 = _zz_currentValidCount_2;
      3'b011 : _zz_currentValidCount_8 = _zz_currentValidCount_3;
      3'b100 : _zz_currentValidCount_8 = _zz_currentValidCount_4;
      3'b101 : _zz_currentValidCount_8 = _zz_currentValidCount_5;
      3'b110 : _zz_currentValidCount_8 = _zz_currentValidCount_6;
      default : _zz_currentValidCount_8 = _zz_currentValidCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_currentValidCount_11)
      3'b000 : _zz_currentValidCount_10 = _zz_currentValidCount;
      3'b001 : _zz_currentValidCount_10 = _zz_currentValidCount_1;
      3'b010 : _zz_currentValidCount_10 = _zz_currentValidCount_2;
      3'b011 : _zz_currentValidCount_10 = _zz_currentValidCount_3;
      3'b100 : _zz_currentValidCount_10 = _zz_currentValidCount_4;
      3'b101 : _zz_currentValidCount_10 = _zz_currentValidCount_5;
      3'b110 : _zz_currentValidCount_10 = _zz_currentValidCount_6;
      default : _zz_currentValidCount_10 = _zz_currentValidCount_7;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : io_allocateIn_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_allocateIn_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_allocateIn_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_allocateIn_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_allocateIn_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_allocateIn_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_allocateIn_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_allocateIn_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_allocateIn_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_allocateIn_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_allocateIn_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_allocateIn_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_allocateIn_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_allocateIn_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_allocateIn_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_allocateIn_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_allocateIn_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_allocateIn_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_allocateIn_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : io_allocateIn_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : io_allocateIn_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_allocateIn_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_allocateIn_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_allocateIn_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_allocateIn_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_allocateIn_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_allocateIn_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_allocateIn_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_isa)
      IsaType_UNKNOWN : io_allocateIn_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_allocateIn_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : io_allocateIn_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_allocateIn_payload_uop_decoded_isa_string = "LOONGARCH";
      default : io_allocateIn_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : io_allocateIn_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_allocateIn_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_allocateIn_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : io_allocateIn_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : io_allocateIn_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "D";
      default : io_allocateIn_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_allocateIn_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_allocateIn_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : io_allocateIn_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocateIn_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : io_allocateIn_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_aluCtrl_logicOp)
      LogicOp_NONE : io_issueOut_payload_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_issueOut_payload_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_issueOut_payload_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_issueOut_payload_aluCtrl_logicOp_string = "XOR_1";
      default : io_issueOut_payload_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_issueOut_payload_immUsage)
      ImmUsageType_NONE : io_issueOut_payload_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_issueOut_payload_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_issueOut_payload_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_issueOut_payload_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_issueOut_payload_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_issueOut_payload_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_issueOut_payload_immUsage_string = "JUMP_OFFSET  ";
      default : io_issueOut_payload_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entries_0_aluCtrl_logicOp)
      LogicOp_NONE : entries_0_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entries_0_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entries_0_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entries_0_aluCtrl_logicOp_string = "XOR_1";
      default : entries_0_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_0_immUsage)
      ImmUsageType_NONE : entries_0_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entries_0_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entries_0_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entries_0_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entries_0_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entries_0_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entries_0_immUsage_string = "JUMP_OFFSET  ";
      default : entries_0_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entries_1_aluCtrl_logicOp)
      LogicOp_NONE : entries_1_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entries_1_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entries_1_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entries_1_aluCtrl_logicOp_string = "XOR_1";
      default : entries_1_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_1_immUsage)
      ImmUsageType_NONE : entries_1_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entries_1_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entries_1_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entries_1_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entries_1_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entries_1_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entries_1_immUsage_string = "JUMP_OFFSET  ";
      default : entries_1_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entries_2_aluCtrl_logicOp)
      LogicOp_NONE : entries_2_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entries_2_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entries_2_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entries_2_aluCtrl_logicOp_string = "XOR_1";
      default : entries_2_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_2_immUsage)
      ImmUsageType_NONE : entries_2_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entries_2_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entries_2_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entries_2_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entries_2_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entries_2_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entries_2_immUsage_string = "JUMP_OFFSET  ";
      default : entries_2_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entries_3_aluCtrl_logicOp)
      LogicOp_NONE : entries_3_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entries_3_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entries_3_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entries_3_aluCtrl_logicOp_string = "XOR_1";
      default : entries_3_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entries_3_immUsage)
      ImmUsageType_NONE : entries_3_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entries_3_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entries_3_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entries_3_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entries_3_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entries_3_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entries_3_immUsage_string = "JUMP_OFFSET  ";
      default : entries_3_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_aluCtrl_logicOp)
      LogicOp_NONE : _zz_io_issueOut_payload_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : _zz_io_issueOut_payload_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : _zz_io_issueOut_payload_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_io_issueOut_payload_aluCtrl_logicOp_string = "XOR_1";
      default : _zz_io_issueOut_payload_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_issueOut_payload_immUsage)
      ImmUsageType_NONE : _zz_io_issueOut_payload_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_io_issueOut_payload_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_io_issueOut_payload_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_io_issueOut_payload_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_io_issueOut_payload_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_io_issueOut_payload_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_io_issueOut_payload_immUsage_string = "JUMP_OFFSET  ";
      default : _zz_io_issueOut_payload_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_aluCtrl_logicOp)
      LogicOp_NONE : entriesNext_0_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entriesNext_0_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entriesNext_0_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entriesNext_0_aluCtrl_logicOp_string = "XOR_1";
      default : entriesNext_0_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_0_immUsage)
      ImmUsageType_NONE : entriesNext_0_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entriesNext_0_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entriesNext_0_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entriesNext_0_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entriesNext_0_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entriesNext_0_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entriesNext_0_immUsage_string = "JUMP_OFFSET  ";
      default : entriesNext_0_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_aluCtrl_logicOp)
      LogicOp_NONE : entriesNext_1_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entriesNext_1_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entriesNext_1_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entriesNext_1_aluCtrl_logicOp_string = "XOR_1";
      default : entriesNext_1_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_1_immUsage)
      ImmUsageType_NONE : entriesNext_1_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entriesNext_1_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entriesNext_1_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entriesNext_1_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entriesNext_1_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entriesNext_1_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entriesNext_1_immUsage_string = "JUMP_OFFSET  ";
      default : entriesNext_1_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_aluCtrl_logicOp)
      LogicOp_NONE : entriesNext_2_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entriesNext_2_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entriesNext_2_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entriesNext_2_aluCtrl_logicOp_string = "XOR_1";
      default : entriesNext_2_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_2_immUsage)
      ImmUsageType_NONE : entriesNext_2_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entriesNext_2_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entriesNext_2_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entriesNext_2_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entriesNext_2_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entriesNext_2_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entriesNext_2_immUsage_string = "JUMP_OFFSET  ";
      default : entriesNext_2_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_aluCtrl_logicOp)
      LogicOp_NONE : entriesNext_3_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : entriesNext_3_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : entriesNext_3_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : entriesNext_3_aluCtrl_logicOp_string = "XOR_1";
      default : entriesNext_3_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(entriesNext_3_immUsage)
      ImmUsageType_NONE : entriesNext_3_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : entriesNext_3_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : entriesNext_3_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : entriesNext_3_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : entriesNext_3_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : entriesNext_3_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : entriesNext_3_immUsage_string = "JUMP_OFFSET  ";
      default : entriesNext_3_immUsage_string = "?????????????";
    endcase
  end
  `endif

  assign io_issueOut_fire = (io_issueOut_valid && io_issueOut_ready);
  assign localWakeupValid = (io_issueOut_fire && io_issueOut_payload_writesToPhysReg);
  always @(*) begin
    wokeUpSrc1Mask = 4'b0000;
    if(entryValids_0) begin
      if(when_IssueQueueComponent_l103) begin
        wokeUpSrc1Mask[0] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_1) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_2) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_3) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_4) begin
          wokeUpSrc1Mask[0] = 1'b1;
        end
      end
    end
    if(entryValids_1) begin
      if(when_IssueQueueComponent_l103_1) begin
        wokeUpSrc1Mask[1] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_5) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_6) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_7) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_8) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_9) begin
          wokeUpSrc1Mask[1] = 1'b1;
        end
      end
    end
    if(entryValids_2) begin
      if(when_IssueQueueComponent_l103_2) begin
        wokeUpSrc1Mask[2] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_10) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_11) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_12) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_13) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_14) begin
          wokeUpSrc1Mask[2] = 1'b1;
        end
      end
    end
    if(entryValids_3) begin
      if(when_IssueQueueComponent_l103_3) begin
        wokeUpSrc1Mask[3] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l113_15) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l113_16) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l113_17) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l113_18) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l113_19) begin
          wokeUpSrc1Mask[3] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    wokeUpSrc2Mask = 4'b0000;
    if(entryValids_0) begin
      if(when_IssueQueueComponent_l106) begin
        wokeUpSrc2Mask[0] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_1) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_2) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_3) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_4) begin
          wokeUpSrc2Mask[0] = 1'b1;
        end
      end
    end
    if(entryValids_1) begin
      if(when_IssueQueueComponent_l106_1) begin
        wokeUpSrc2Mask[1] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_5) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_6) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_7) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_8) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_9) begin
          wokeUpSrc2Mask[1] = 1'b1;
        end
      end
    end
    if(entryValids_2) begin
      if(when_IssueQueueComponent_l106_2) begin
        wokeUpSrc2Mask[2] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_10) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_11) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_12) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_13) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_14) begin
          wokeUpSrc2Mask[2] = 1'b1;
        end
      end
    end
    if(entryValids_3) begin
      if(when_IssueQueueComponent_l106_3) begin
        wokeUpSrc2Mask[3] = 1'b1;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l116_15) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l116_16) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l116_17) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l116_18) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l116_19) begin
          wokeUpSrc2Mask[3] = 1'b1;
        end
      end
    end
  end

  assign _zz_when_IssueQueueComponent_l103 = ((! entries_0_src1Ready) && entries_0_useSrc1);
  assign _zz_when_IssueQueueComponent_l106 = ((! entries_0_src2Ready) && entries_0_useSrc2);
  assign when_IssueQueueComponent_l103 = ((_zz_when_IssueQueueComponent_l103 && localWakeupValid) && (entries_0_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106 = ((_zz_when_IssueQueueComponent_l106 && localWakeupValid) && (entries_0_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_1 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_1 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_2 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_2 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_3 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_3 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_4 = (_zz_when_IssueQueueComponent_l103 && (entries_0_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_4 = (_zz_when_IssueQueueComponent_l106 && (entries_0_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_1 = ((! entries_1_src1Ready) && entries_1_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_1 = ((! entries_1_src2Ready) && entries_1_useSrc2);
  assign when_IssueQueueComponent_l103_1 = ((_zz_when_IssueQueueComponent_l103_1 && localWakeupValid) && (entries_1_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_1 = ((_zz_when_IssueQueueComponent_l106_1 && localWakeupValid) && (entries_1_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_5 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_5 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_6 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_6 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_7 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_7 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_8 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_8 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_9 = (_zz_when_IssueQueueComponent_l103_1 && (entries_1_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_9 = (_zz_when_IssueQueueComponent_l106_1 && (entries_1_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_2 = ((! entries_2_src1Ready) && entries_2_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_2 = ((! entries_2_src2Ready) && entries_2_useSrc2);
  assign when_IssueQueueComponent_l103_2 = ((_zz_when_IssueQueueComponent_l103_2 && localWakeupValid) && (entries_2_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_2 = ((_zz_when_IssueQueueComponent_l106_2 && localWakeupValid) && (entries_2_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_10 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_10 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_11 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_11 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_12 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_12 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_13 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_13 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_14 = (_zz_when_IssueQueueComponent_l103_2 && (entries_2_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_14 = (_zz_when_IssueQueueComponent_l106_2 && (entries_2_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_when_IssueQueueComponent_l103_3 = ((! entries_3_src1Ready) && entries_3_useSrc1);
  assign _zz_when_IssueQueueComponent_l106_3 = ((! entries_3_src2Ready) && entries_3_useSrc2);
  assign when_IssueQueueComponent_l103_3 = ((_zz_when_IssueQueueComponent_l103_3 && localWakeupValid) && (entries_3_src1Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l106_3 = ((_zz_when_IssueQueueComponent_l106_3 && localWakeupValid) && (entries_3_src2Tag == io_issueOut_payload_physDest_idx));
  assign when_IssueQueueComponent_l113_15 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_15 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_16 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_16 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_17 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_17 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_18 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_18 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l113_19 = (_zz_when_IssueQueueComponent_l103_3 && (entries_3_src1Tag == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l116_19 = (_zz_when_IssueQueueComponent_l106_3 && (entries_3_src2Tag == io_wakeupIn_4_payload_physRegIdx));
  assign entriesReadyToIssue_0 = ((entryValids_0 && ((! entries_0_useSrc1) || entries_0_src1Ready)) && ((! entries_0_useSrc2) || entries_0_src2Ready));
  assign entriesReadyToIssue_1 = ((entryValids_1 && ((! entries_1_useSrc1) || entries_1_src1Ready)) && ((! entries_1_useSrc2) || entries_1_src2Ready));
  assign entriesReadyToIssue_2 = ((entryValids_2 && ((! entries_2_useSrc1) || entries_2_src1Ready)) && ((! entries_2_useSrc2) || entries_2_src2Ready));
  assign entriesReadyToIssue_3 = ((entryValids_3 && ((! entries_3_useSrc1) || entries_3_src1Ready)) && ((! entries_3_useSrc2) || entries_3_src2Ready));
  assign issueRequestMask = {entriesReadyToIssue_3,{entriesReadyToIssue_2,{entriesReadyToIssue_1,entriesReadyToIssue_0}}};
  assign issueRequestMask_ohFirst_input = issueRequestMask;
  assign issueRequestMask_ohFirst_masked = (issueRequestMask_ohFirst_input & (~ _zz_issueRequestMask_ohFirst_masked));
  assign issueRequestOh = issueRequestMask_ohFirst_masked;
  assign _zz_issueIdx = issueRequestOh[3];
  assign _zz_issueIdx_1 = (issueRequestOh[1] || _zz_issueIdx);
  assign _zz_issueIdx_2 = (issueRequestOh[2] || _zz_issueIdx);
  assign issueIdx = {_zz_issueIdx_2,_zz_issueIdx_1};
  assign io_issueOut_valid = ((|issueRequestOh) && (! io_flush));
  assign _zz_io_issueOut_payload_aluCtrl_logicOp = _zz__zz_io_issueOut_payload_aluCtrl_logicOp;
  assign _zz_io_issueOut_payload_immUsage = _zz__zz_io_issueOut_payload_immUsage;
  assign io_issueOut_payload_robPtr = _zz_io_issueOut_payload_robPtr;
  assign io_issueOut_payload_physDest_idx = _zz_io_issueOut_payload_physDest_idx;
  assign io_issueOut_payload_physDestIsFpr = _zz_io_issueOut_payload_physDestIsFpr;
  assign io_issueOut_payload_writesToPhysReg = _zz_io_issueOut_payload_writesToPhysReg;
  assign io_issueOut_payload_useSrc1 = _zz_io_issueOut_payload_useSrc1;
  assign io_issueOut_payload_src1Data = _zz_io_issueOut_payload_src1Data;
  assign io_issueOut_payload_src1Tag = _zz_io_issueOut_payload_src1Tag;
  assign io_issueOut_payload_src1Ready = _zz_io_issueOut_payload_src1Ready;
  assign io_issueOut_payload_src1IsFpr = _zz_io_issueOut_payload_src1IsFpr;
  assign io_issueOut_payload_useSrc2 = _zz_io_issueOut_payload_useSrc2;
  assign io_issueOut_payload_src2Data = _zz_io_issueOut_payload_src2Data;
  assign io_issueOut_payload_src2Tag = _zz_io_issueOut_payload_src2Tag;
  assign io_issueOut_payload_src2Ready = _zz_io_issueOut_payload_src2Ready;
  assign io_issueOut_payload_src2IsFpr = _zz_io_issueOut_payload_src2IsFpr;
  assign io_issueOut_payload_aluCtrl_valid = _zz_io_issueOut_payload_aluCtrl_valid;
  assign io_issueOut_payload_aluCtrl_isSub = _zz_io_issueOut_payload_aluCtrl_isSub;
  assign io_issueOut_payload_aluCtrl_isAdd = _zz_io_issueOut_payload_aluCtrl_isAdd;
  assign io_issueOut_payload_aluCtrl_isSigned = _zz_io_issueOut_payload_aluCtrl_isSigned;
  assign io_issueOut_payload_aluCtrl_logicOp = _zz_io_issueOut_payload_aluCtrl_logicOp;
  assign io_issueOut_payload_shiftCtrl_valid = _zz_io_issueOut_payload_shiftCtrl_valid;
  assign io_issueOut_payload_shiftCtrl_isRight = _zz_io_issueOut_payload_shiftCtrl_isRight;
  assign io_issueOut_payload_shiftCtrl_isArithmetic = _zz_io_issueOut_payload_shiftCtrl_isArithmetic;
  assign io_issueOut_payload_shiftCtrl_isRotate = _zz_io_issueOut_payload_shiftCtrl_isRotate;
  assign io_issueOut_payload_shiftCtrl_isDoubleWord = _zz_io_issueOut_payload_shiftCtrl_isDoubleWord;
  assign io_issueOut_payload_imm = _zz_io_issueOut_payload_imm;
  assign io_issueOut_payload_immUsage = _zz_io_issueOut_payload_immUsage;
  assign freeSlotsMask = {(! entryValids_3),{(! entryValids_2),{(! entryValids_1),(! entryValids_0)}}};
  assign hasSpaceForNewEntry = ((|freeSlotsMask) || io_issueOut_fire);
  assign io_allocateIn_ready = (hasSpaceForNewEntry && (! io_flush));
  always @(*) begin
    firedSlotMask = 4'b0000;
    if(io_issueOut_fire) begin
      firedSlotMask[issueIdx] = 1'b1;
    end
  end

  assign _zz_allocationMask = (freeSlotsMask | firedSlotMask);
  assign allocationMask = (_zz_allocationMask & (~ _zz_allocationMask_1));
  assign _zz_allocateIdx = allocationMask[3];
  assign _zz_allocateIdx_1 = (allocationMask[1] || _zz_allocateIdx);
  assign _zz_allocateIdx_2 = (allocationMask[2] || _zz_allocateIdx);
  assign allocateIdx = {_zz_allocateIdx_2,_zz_allocateIdx_1};
  always @(*) begin
    entriesNext_0_robPtr = entries_0_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_physDest_idx = entries_0_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_physDestIsFpr = entries_0_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_writesToPhysReg = entries_0_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_0_useSrc1 = entries_0_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Data = entries_0_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Tag = entries_0_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1Ready = entries_0_src1Ready;
    if(when_IssueQueueComponent_l186) begin
      entriesNext_0_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_3) begin
        entriesNext_0_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_3) begin
            entriesNext_0_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_0_src1IsFpr = entries_0_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_useSrc2 = entries_0_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Data = entries_0_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Tag = entries_0_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2Ready = entries_0_src2Ready;
    if(when_IssueQueueComponent_l187) begin
      entriesNext_0_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_3) begin
        entriesNext_0_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_3) begin
            entriesNext_0_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_0_src2IsFpr = entries_0_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_0_aluCtrl_valid = entries_0_aluCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_aluCtrl_valid = io_allocateIn_payload_uop_decoded_aluCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_0_aluCtrl_isSub = entries_0_aluCtrl_isSub;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_aluCtrl_isSub = io_allocateIn_payload_uop_decoded_aluCtrl_isSub;
      end
    end
  end

  always @(*) begin
    entriesNext_0_aluCtrl_isAdd = entries_0_aluCtrl_isAdd;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_aluCtrl_isAdd = io_allocateIn_payload_uop_decoded_aluCtrl_isAdd;
      end
    end
  end

  always @(*) begin
    entriesNext_0_aluCtrl_isSigned = entries_0_aluCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_aluCtrl_isSigned = io_allocateIn_payload_uop_decoded_aluCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_0_aluCtrl_logicOp = entries_0_aluCtrl_logicOp;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_aluCtrl_logicOp = io_allocateIn_payload_uop_decoded_aluCtrl_logicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_0_shiftCtrl_valid = entries_0_shiftCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_shiftCtrl_valid = io_allocateIn_payload_uop_decoded_shiftCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_0_shiftCtrl_isRight = entries_0_shiftCtrl_isRight;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_shiftCtrl_isRight = io_allocateIn_payload_uop_decoded_shiftCtrl_isRight;
      end
    end
  end

  always @(*) begin
    entriesNext_0_shiftCtrl_isArithmetic = entries_0_shiftCtrl_isArithmetic;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_shiftCtrl_isArithmetic = io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic;
      end
    end
  end

  always @(*) begin
    entriesNext_0_shiftCtrl_isRotate = entries_0_shiftCtrl_isRotate;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_shiftCtrl_isRotate = io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate;
      end
    end
  end

  always @(*) begin
    entriesNext_0_shiftCtrl_isDoubleWord = entries_0_shiftCtrl_isDoubleWord;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_shiftCtrl_isDoubleWord = io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord;
      end
    end
  end

  always @(*) begin
    entriesNext_0_imm = entries_0_imm;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_0_immUsage = entries_0_immUsage;
    if(io_allocateIn_fire) begin
      if(_zz_3) begin
        entriesNext_0_immUsage = io_allocateIn_payload_uop_decoded_immUsage;
      end
    end
  end

  always @(*) begin
    entriesNext_1_robPtr = entries_1_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_physDest_idx = entries_1_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_physDestIsFpr = entries_1_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_writesToPhysReg = entries_1_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_1_useSrc1 = entries_1_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Data = entries_1_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Tag = entries_1_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1Ready = entries_1_src1Ready;
    if(when_IssueQueueComponent_l186_1) begin
      entriesNext_1_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_4) begin
        entriesNext_1_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_4) begin
            entriesNext_1_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_1_src1IsFpr = entries_1_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_useSrc2 = entries_1_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Data = entries_1_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Tag = entries_1_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2Ready = entries_1_src2Ready;
    if(when_IssueQueueComponent_l187_1) begin
      entriesNext_1_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_4) begin
        entriesNext_1_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_4) begin
            entriesNext_1_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_1_src2IsFpr = entries_1_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_1_aluCtrl_valid = entries_1_aluCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_aluCtrl_valid = io_allocateIn_payload_uop_decoded_aluCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_1_aluCtrl_isSub = entries_1_aluCtrl_isSub;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_aluCtrl_isSub = io_allocateIn_payload_uop_decoded_aluCtrl_isSub;
      end
    end
  end

  always @(*) begin
    entriesNext_1_aluCtrl_isAdd = entries_1_aluCtrl_isAdd;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_aluCtrl_isAdd = io_allocateIn_payload_uop_decoded_aluCtrl_isAdd;
      end
    end
  end

  always @(*) begin
    entriesNext_1_aluCtrl_isSigned = entries_1_aluCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_aluCtrl_isSigned = io_allocateIn_payload_uop_decoded_aluCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_1_aluCtrl_logicOp = entries_1_aluCtrl_logicOp;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_aluCtrl_logicOp = io_allocateIn_payload_uop_decoded_aluCtrl_logicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_1_shiftCtrl_valid = entries_1_shiftCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_shiftCtrl_valid = io_allocateIn_payload_uop_decoded_shiftCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_1_shiftCtrl_isRight = entries_1_shiftCtrl_isRight;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_shiftCtrl_isRight = io_allocateIn_payload_uop_decoded_shiftCtrl_isRight;
      end
    end
  end

  always @(*) begin
    entriesNext_1_shiftCtrl_isArithmetic = entries_1_shiftCtrl_isArithmetic;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_shiftCtrl_isArithmetic = io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic;
      end
    end
  end

  always @(*) begin
    entriesNext_1_shiftCtrl_isRotate = entries_1_shiftCtrl_isRotate;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_shiftCtrl_isRotate = io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate;
      end
    end
  end

  always @(*) begin
    entriesNext_1_shiftCtrl_isDoubleWord = entries_1_shiftCtrl_isDoubleWord;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_shiftCtrl_isDoubleWord = io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord;
      end
    end
  end

  always @(*) begin
    entriesNext_1_imm = entries_1_imm;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_1_immUsage = entries_1_immUsage;
    if(io_allocateIn_fire) begin
      if(_zz_4) begin
        entriesNext_1_immUsage = io_allocateIn_payload_uop_decoded_immUsage;
      end
    end
  end

  always @(*) begin
    entriesNext_2_robPtr = entries_2_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_physDest_idx = entries_2_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_physDestIsFpr = entries_2_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_writesToPhysReg = entries_2_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_2_useSrc1 = entries_2_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Data = entries_2_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Tag = entries_2_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1Ready = entries_2_src1Ready;
    if(when_IssueQueueComponent_l186_2) begin
      entriesNext_2_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_5) begin
        entriesNext_2_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_5) begin
            entriesNext_2_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_2_src1IsFpr = entries_2_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_useSrc2 = entries_2_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Data = entries_2_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Tag = entries_2_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2Ready = entries_2_src2Ready;
    if(when_IssueQueueComponent_l187_2) begin
      entriesNext_2_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_5) begin
        entriesNext_2_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_5) begin
            entriesNext_2_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_2_src2IsFpr = entries_2_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_2_aluCtrl_valid = entries_2_aluCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_aluCtrl_valid = io_allocateIn_payload_uop_decoded_aluCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_2_aluCtrl_isSub = entries_2_aluCtrl_isSub;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_aluCtrl_isSub = io_allocateIn_payload_uop_decoded_aluCtrl_isSub;
      end
    end
  end

  always @(*) begin
    entriesNext_2_aluCtrl_isAdd = entries_2_aluCtrl_isAdd;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_aluCtrl_isAdd = io_allocateIn_payload_uop_decoded_aluCtrl_isAdd;
      end
    end
  end

  always @(*) begin
    entriesNext_2_aluCtrl_isSigned = entries_2_aluCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_aluCtrl_isSigned = io_allocateIn_payload_uop_decoded_aluCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_2_aluCtrl_logicOp = entries_2_aluCtrl_logicOp;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_aluCtrl_logicOp = io_allocateIn_payload_uop_decoded_aluCtrl_logicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_2_shiftCtrl_valid = entries_2_shiftCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_shiftCtrl_valid = io_allocateIn_payload_uop_decoded_shiftCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_2_shiftCtrl_isRight = entries_2_shiftCtrl_isRight;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_shiftCtrl_isRight = io_allocateIn_payload_uop_decoded_shiftCtrl_isRight;
      end
    end
  end

  always @(*) begin
    entriesNext_2_shiftCtrl_isArithmetic = entries_2_shiftCtrl_isArithmetic;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_shiftCtrl_isArithmetic = io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic;
      end
    end
  end

  always @(*) begin
    entriesNext_2_shiftCtrl_isRotate = entries_2_shiftCtrl_isRotate;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_shiftCtrl_isRotate = io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate;
      end
    end
  end

  always @(*) begin
    entriesNext_2_shiftCtrl_isDoubleWord = entries_2_shiftCtrl_isDoubleWord;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_shiftCtrl_isDoubleWord = io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord;
      end
    end
  end

  always @(*) begin
    entriesNext_2_imm = entries_2_imm;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_2_immUsage = entries_2_immUsage;
    if(io_allocateIn_fire) begin
      if(_zz_5) begin
        entriesNext_2_immUsage = io_allocateIn_payload_uop_decoded_immUsage;
      end
    end
  end

  always @(*) begin
    entriesNext_3_robPtr = entries_3_robPtr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_robPtr = io_allocateIn_payload_uop_robPtr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_physDest_idx = entries_3_physDest_idx;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_physDest_idx = io_allocateIn_payload_uop_rename_physDest_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_physDestIsFpr = entries_3_physDestIsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_physDestIsFpr = io_allocateIn_payload_uop_rename_physDestIsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_writesToPhysReg = entries_3_writesToPhysReg;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_writesToPhysReg = io_allocateIn_payload_uop_rename_writesToPhysReg;
      end
    end
  end

  always @(*) begin
    entriesNext_3_useSrc1 = entries_3_useSrc1;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_useSrc1 = io_allocateIn_payload_uop_decoded_useArchSrc1;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Data = entries_3_src1Data;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Tag = entries_3_src1Tag;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Tag = io_allocateIn_payload_uop_rename_physSrc1_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1Ready = entries_3_src1Ready;
    if(when_IssueQueueComponent_l186_3) begin
      entriesNext_3_src1Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1Ready = _zz_entriesNext_0_src1Ready;
      end
      if(_zz_6) begin
        entriesNext_3_src1Ready = io_allocateIn_payload_src1InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l212) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l212_1) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l212_2) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l212_3) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l212_4) begin
          if(_zz_6) begin
            entriesNext_3_src1Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_3_src1IsFpr = entries_3_src1IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src1IsFpr = io_allocateIn_payload_uop_rename_physSrc1IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_useSrc2 = entries_3_useSrc2;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_useSrc2 = io_allocateIn_payload_uop_decoded_useArchSrc2;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Data = entries_3_src2Data;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Tag = entries_3_src2Tag;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Tag = io_allocateIn_payload_uop_rename_physSrc2_idx;
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2Ready = entries_3_src2Ready;
    if(when_IssueQueueComponent_l187_3) begin
      entriesNext_3_src2Ready = 1'b1;
    end
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2Ready = _zz_entriesNext_0_src2Ready;
      end
      if(_zz_6) begin
        entriesNext_3_src2Ready = io_allocateIn_payload_src2InitialReady;
      end
      if(io_wakeupIn_0_valid) begin
        if(when_IssueQueueComponent_l215) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_1_valid) begin
        if(when_IssueQueueComponent_l215_1) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_2_valid) begin
        if(when_IssueQueueComponent_l215_2) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_3_valid) begin
        if(when_IssueQueueComponent_l215_3) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
      if(io_wakeupIn_4_valid) begin
        if(when_IssueQueueComponent_l215_4) begin
          if(_zz_6) begin
            entriesNext_3_src2Ready = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    entriesNext_3_src2IsFpr = entries_3_src2IsFpr;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_src2IsFpr = io_allocateIn_payload_uop_rename_physSrc2IsFpr;
      end
    end
  end

  always @(*) begin
    entriesNext_3_aluCtrl_valid = entries_3_aluCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_aluCtrl_valid = io_allocateIn_payload_uop_decoded_aluCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_3_aluCtrl_isSub = entries_3_aluCtrl_isSub;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_aluCtrl_isSub = io_allocateIn_payload_uop_decoded_aluCtrl_isSub;
      end
    end
  end

  always @(*) begin
    entriesNext_3_aluCtrl_isAdd = entries_3_aluCtrl_isAdd;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_aluCtrl_isAdd = io_allocateIn_payload_uop_decoded_aluCtrl_isAdd;
      end
    end
  end

  always @(*) begin
    entriesNext_3_aluCtrl_isSigned = entries_3_aluCtrl_isSigned;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_aluCtrl_isSigned = io_allocateIn_payload_uop_decoded_aluCtrl_isSigned;
      end
    end
  end

  always @(*) begin
    entriesNext_3_aluCtrl_logicOp = entries_3_aluCtrl_logicOp;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_aluCtrl_logicOp = io_allocateIn_payload_uop_decoded_aluCtrl_logicOp;
      end
    end
  end

  always @(*) begin
    entriesNext_3_shiftCtrl_valid = entries_3_shiftCtrl_valid;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_shiftCtrl_valid = io_allocateIn_payload_uop_decoded_shiftCtrl_valid;
      end
    end
  end

  always @(*) begin
    entriesNext_3_shiftCtrl_isRight = entries_3_shiftCtrl_isRight;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_shiftCtrl_isRight = io_allocateIn_payload_uop_decoded_shiftCtrl_isRight;
      end
    end
  end

  always @(*) begin
    entriesNext_3_shiftCtrl_isArithmetic = entries_3_shiftCtrl_isArithmetic;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_shiftCtrl_isArithmetic = io_allocateIn_payload_uop_decoded_shiftCtrl_isArithmetic;
      end
    end
  end

  always @(*) begin
    entriesNext_3_shiftCtrl_isRotate = entries_3_shiftCtrl_isRotate;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_shiftCtrl_isRotate = io_allocateIn_payload_uop_decoded_shiftCtrl_isRotate;
      end
    end
  end

  always @(*) begin
    entriesNext_3_shiftCtrl_isDoubleWord = entries_3_shiftCtrl_isDoubleWord;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_shiftCtrl_isDoubleWord = io_allocateIn_payload_uop_decoded_shiftCtrl_isDoubleWord;
      end
    end
  end

  always @(*) begin
    entriesNext_3_imm = entries_3_imm;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_imm = io_allocateIn_payload_uop_decoded_imm;
      end
    end
  end

  always @(*) begin
    entriesNext_3_immUsage = entries_3_immUsage;
    if(io_allocateIn_fire) begin
      if(_zz_6) begin
        entriesNext_3_immUsage = io_allocateIn_payload_uop_decoded_immUsage;
      end
    end
  end

  always @(*) begin
    entryValidsNext_0 = entryValids_0;
    if(io_issueOut_fire) begin
      if(_zz_1[0]) begin
        entryValidsNext_0 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[0]) begin
        entryValidsNext_0 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_0 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_1 = entryValids_1;
    if(io_issueOut_fire) begin
      if(_zz_1[1]) begin
        entryValidsNext_1 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[1]) begin
        entryValidsNext_1 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_1 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_2 = entryValids_2;
    if(io_issueOut_fire) begin
      if(_zz_1[2]) begin
        entryValidsNext_2 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[2]) begin
        entryValidsNext_2 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_2 = 1'b0;
    end
  end

  always @(*) begin
    entryValidsNext_3 = entryValids_3;
    if(io_issueOut_fire) begin
      if(_zz_1[3]) begin
        entryValidsNext_3 = 1'b0;
      end
    end
    if(io_allocateIn_fire) begin
      if(_zz_7[3]) begin
        entryValidsNext_3 = 1'b1;
      end
    end
    if(io_flush) begin
      entryValidsNext_3 = 1'b0;
    end
  end

  assign when_IssueQueueComponent_l186 = wokeUpSrc1Mask[0];
  assign when_IssueQueueComponent_l187 = wokeUpSrc2Mask[0];
  assign when_IssueQueueComponent_l186_1 = wokeUpSrc1Mask[1];
  assign when_IssueQueueComponent_l187_1 = wokeUpSrc2Mask[1];
  assign when_IssueQueueComponent_l186_2 = wokeUpSrc1Mask[2];
  assign when_IssueQueueComponent_l187_2 = wokeUpSrc2Mask[2];
  assign when_IssueQueueComponent_l186_3 = wokeUpSrc1Mask[3];
  assign when_IssueQueueComponent_l187_3 = wokeUpSrc2Mask[3];
  assign _zz_1 = ({3'd0,1'b1} <<< issueIdx);
  assign io_allocateIn_fire = (io_allocateIn_valid && io_allocateIn_ready);
  assign _zz_2 = ({3'd0,1'b1} <<< allocateIdx);
  assign _zz_3 = _zz_2[0];
  assign _zz_4 = _zz_2[1];
  assign _zz_5 = _zz_2[2];
  assign _zz_6 = _zz_2[3];
  assign _zz_entriesNext_0_src1Ready = (! io_allocateIn_payload_uop_decoded_useArchSrc1);
  assign _zz_entriesNext_0_src2Ready = (! io_allocateIn_payload_uop_decoded_useArchSrc2);
  assign _zz_7 = ({3'd0,1'b1} <<< allocateIdx);
  assign when_IssueQueueComponent_l212 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l215 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_0_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_1 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_1 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_1_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_2 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_2 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_2_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_3 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_3 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_3_payload_physRegIdx));
  assign when_IssueQueueComponent_l212_4 = ((io_allocateIn_payload_uop_decoded_useArchSrc1 && (! io_allocateIn_payload_src1InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc1_idx == io_wakeupIn_4_payload_physRegIdx));
  assign when_IssueQueueComponent_l215_4 = ((io_allocateIn_payload_uop_decoded_useArchSrc2 && (! io_allocateIn_payload_src2InitialReady)) && (io_allocateIn_payload_uop_rename_physSrc2_idx == io_wakeupIn_4_payload_physRegIdx));
  assign _zz_currentValidCount = 3'b000;
  assign _zz_currentValidCount_1 = 3'b001;
  assign _zz_currentValidCount_2 = 3'b001;
  assign _zz_currentValidCount_3 = 3'b010;
  assign _zz_currentValidCount_4 = 3'b001;
  assign _zz_currentValidCount_5 = 3'b010;
  assign _zz_currentValidCount_6 = 3'b010;
  assign _zz_currentValidCount_7 = 3'b011;
  assign currentValidCount = (_zz_currentValidCount_8 + _zz_currentValidCount_10);
  assign logCondition = (io_allocateIn_fire || io_issueOut_fire);
  assign when_IssueQueueComponent_l256 = (logCondition && (3'b000 < currentValidCount));
  always @(posedge clk) begin
    if(reset) begin
      entryValids_0 <= 1'b0;
      entryValids_1 <= 1'b0;
      entryValids_2 <= 1'b0;
      entryValids_3 <= 1'b0;
    end else begin
      entryValids_0 <= entryValidsNext_0;
      entryValids_1 <= entryValidsNext_1;
      entryValids_2 <= entryValidsNext_2;
      entryValids_3 <= entryValidsNext_3;
      if(logCondition) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // IssueQueueComponent.scala:L247
          `else
            if(!1'b0) begin
              $display("NOTE(IssueQueueComponent.scala:247):  [normal] AluIntEU_IQ-0: STATUS - ValidCount=%x, allocateIn(valid=%x, ready=%x), issueOut(valid=%x, ready=%x)", currentValidCount, io_allocateIn_valid, io_allocateIn_ready, io_issueOut_valid, io_issueOut_ready); // IssueQueueComponent.scala:L247
            end
          `endif
        `endif
      end
      if(when_IssueQueueComponent_l256) begin
        if(entryValids_0) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] AluIntEU_IQ-0: (LAST CYCLE) ENTRY[0] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_0_robPtr, entries_0_physDest_idx, entries_0_useSrc1, entries_0_src1Tag, entries_0_src1Ready, entries_0_useSrc2, entries_0_src2Tag, entries_0_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_1) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] AluIntEU_IQ-0: (LAST CYCLE) ENTRY[1] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_1_robPtr, entries_1_physDest_idx, entries_1_useSrc1, entries_1_src1Tag, entries_1_src1Ready, entries_1_useSrc2, entries_1_src2Tag, entries_1_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_2) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] AluIntEU_IQ-0: (LAST CYCLE) ENTRY[2] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_2_robPtr, entries_2_physDest_idx, entries_2_useSrc1, entries_2_src1Tag, entries_2_src1Ready, entries_2_useSrc2, entries_2_src2Tag, entries_2_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
        if(entryValids_3) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // IssueQueueComponent.scala:L259
            `else
              if(!1'b0) begin
                $display("NOTE(IssueQueueComponent.scala:259):  [normal] AluIntEU_IQ-0: (LAST CYCLE) ENTRY[3] - RobPtr=%x, PhysDest=%x, UseSrc1=%x, Src1Tag=%x, Src1Ready=%x, UseSrc2=%x, Src2Tag=%x, Src2Ready=%x", entries_3_robPtr, entries_3_physDest_idx, entries_3_useSrc1, entries_3_src1Tag, entries_3_src1Ready, entries_3_useSrc2, entries_3_src2Tag, entries_3_src2Ready); // IssueQueueComponent.scala:L259
              end
            `endif
          `endif
        end
      end
    end
  end

  always @(posedge clk) begin
    entries_0_robPtr <= entriesNext_0_robPtr;
    entries_0_physDest_idx <= entriesNext_0_physDest_idx;
    entries_0_physDestIsFpr <= entriesNext_0_physDestIsFpr;
    entries_0_writesToPhysReg <= entriesNext_0_writesToPhysReg;
    entries_0_useSrc1 <= entriesNext_0_useSrc1;
    entries_0_src1Data <= entriesNext_0_src1Data;
    entries_0_src1Tag <= entriesNext_0_src1Tag;
    entries_0_src1Ready <= entriesNext_0_src1Ready;
    entries_0_src1IsFpr <= entriesNext_0_src1IsFpr;
    entries_0_useSrc2 <= entriesNext_0_useSrc2;
    entries_0_src2Data <= entriesNext_0_src2Data;
    entries_0_src2Tag <= entriesNext_0_src2Tag;
    entries_0_src2Ready <= entriesNext_0_src2Ready;
    entries_0_src2IsFpr <= entriesNext_0_src2IsFpr;
    entries_0_aluCtrl_valid <= entriesNext_0_aluCtrl_valid;
    entries_0_aluCtrl_isSub <= entriesNext_0_aluCtrl_isSub;
    entries_0_aluCtrl_isAdd <= entriesNext_0_aluCtrl_isAdd;
    entries_0_aluCtrl_isSigned <= entriesNext_0_aluCtrl_isSigned;
    entries_0_aluCtrl_logicOp <= entriesNext_0_aluCtrl_logicOp;
    entries_0_shiftCtrl_valid <= entriesNext_0_shiftCtrl_valid;
    entries_0_shiftCtrl_isRight <= entriesNext_0_shiftCtrl_isRight;
    entries_0_shiftCtrl_isArithmetic <= entriesNext_0_shiftCtrl_isArithmetic;
    entries_0_shiftCtrl_isRotate <= entriesNext_0_shiftCtrl_isRotate;
    entries_0_shiftCtrl_isDoubleWord <= entriesNext_0_shiftCtrl_isDoubleWord;
    entries_0_imm <= entriesNext_0_imm;
    entries_0_immUsage <= entriesNext_0_immUsage;
    entries_1_robPtr <= entriesNext_1_robPtr;
    entries_1_physDest_idx <= entriesNext_1_physDest_idx;
    entries_1_physDestIsFpr <= entriesNext_1_physDestIsFpr;
    entries_1_writesToPhysReg <= entriesNext_1_writesToPhysReg;
    entries_1_useSrc1 <= entriesNext_1_useSrc1;
    entries_1_src1Data <= entriesNext_1_src1Data;
    entries_1_src1Tag <= entriesNext_1_src1Tag;
    entries_1_src1Ready <= entriesNext_1_src1Ready;
    entries_1_src1IsFpr <= entriesNext_1_src1IsFpr;
    entries_1_useSrc2 <= entriesNext_1_useSrc2;
    entries_1_src2Data <= entriesNext_1_src2Data;
    entries_1_src2Tag <= entriesNext_1_src2Tag;
    entries_1_src2Ready <= entriesNext_1_src2Ready;
    entries_1_src2IsFpr <= entriesNext_1_src2IsFpr;
    entries_1_aluCtrl_valid <= entriesNext_1_aluCtrl_valid;
    entries_1_aluCtrl_isSub <= entriesNext_1_aluCtrl_isSub;
    entries_1_aluCtrl_isAdd <= entriesNext_1_aluCtrl_isAdd;
    entries_1_aluCtrl_isSigned <= entriesNext_1_aluCtrl_isSigned;
    entries_1_aluCtrl_logicOp <= entriesNext_1_aluCtrl_logicOp;
    entries_1_shiftCtrl_valid <= entriesNext_1_shiftCtrl_valid;
    entries_1_shiftCtrl_isRight <= entriesNext_1_shiftCtrl_isRight;
    entries_1_shiftCtrl_isArithmetic <= entriesNext_1_shiftCtrl_isArithmetic;
    entries_1_shiftCtrl_isRotate <= entriesNext_1_shiftCtrl_isRotate;
    entries_1_shiftCtrl_isDoubleWord <= entriesNext_1_shiftCtrl_isDoubleWord;
    entries_1_imm <= entriesNext_1_imm;
    entries_1_immUsage <= entriesNext_1_immUsage;
    entries_2_robPtr <= entriesNext_2_robPtr;
    entries_2_physDest_idx <= entriesNext_2_physDest_idx;
    entries_2_physDestIsFpr <= entriesNext_2_physDestIsFpr;
    entries_2_writesToPhysReg <= entriesNext_2_writesToPhysReg;
    entries_2_useSrc1 <= entriesNext_2_useSrc1;
    entries_2_src1Data <= entriesNext_2_src1Data;
    entries_2_src1Tag <= entriesNext_2_src1Tag;
    entries_2_src1Ready <= entriesNext_2_src1Ready;
    entries_2_src1IsFpr <= entriesNext_2_src1IsFpr;
    entries_2_useSrc2 <= entriesNext_2_useSrc2;
    entries_2_src2Data <= entriesNext_2_src2Data;
    entries_2_src2Tag <= entriesNext_2_src2Tag;
    entries_2_src2Ready <= entriesNext_2_src2Ready;
    entries_2_src2IsFpr <= entriesNext_2_src2IsFpr;
    entries_2_aluCtrl_valid <= entriesNext_2_aluCtrl_valid;
    entries_2_aluCtrl_isSub <= entriesNext_2_aluCtrl_isSub;
    entries_2_aluCtrl_isAdd <= entriesNext_2_aluCtrl_isAdd;
    entries_2_aluCtrl_isSigned <= entriesNext_2_aluCtrl_isSigned;
    entries_2_aluCtrl_logicOp <= entriesNext_2_aluCtrl_logicOp;
    entries_2_shiftCtrl_valid <= entriesNext_2_shiftCtrl_valid;
    entries_2_shiftCtrl_isRight <= entriesNext_2_shiftCtrl_isRight;
    entries_2_shiftCtrl_isArithmetic <= entriesNext_2_shiftCtrl_isArithmetic;
    entries_2_shiftCtrl_isRotate <= entriesNext_2_shiftCtrl_isRotate;
    entries_2_shiftCtrl_isDoubleWord <= entriesNext_2_shiftCtrl_isDoubleWord;
    entries_2_imm <= entriesNext_2_imm;
    entries_2_immUsage <= entriesNext_2_immUsage;
    entries_3_robPtr <= entriesNext_3_robPtr;
    entries_3_physDest_idx <= entriesNext_3_physDest_idx;
    entries_3_physDestIsFpr <= entriesNext_3_physDestIsFpr;
    entries_3_writesToPhysReg <= entriesNext_3_writesToPhysReg;
    entries_3_useSrc1 <= entriesNext_3_useSrc1;
    entries_3_src1Data <= entriesNext_3_src1Data;
    entries_3_src1Tag <= entriesNext_3_src1Tag;
    entries_3_src1Ready <= entriesNext_3_src1Ready;
    entries_3_src1IsFpr <= entriesNext_3_src1IsFpr;
    entries_3_useSrc2 <= entriesNext_3_useSrc2;
    entries_3_src2Data <= entriesNext_3_src2Data;
    entries_3_src2Tag <= entriesNext_3_src2Tag;
    entries_3_src2Ready <= entriesNext_3_src2Ready;
    entries_3_src2IsFpr <= entriesNext_3_src2IsFpr;
    entries_3_aluCtrl_valid <= entriesNext_3_aluCtrl_valid;
    entries_3_aluCtrl_isSub <= entriesNext_3_aluCtrl_isSub;
    entries_3_aluCtrl_isAdd <= entriesNext_3_aluCtrl_isAdd;
    entries_3_aluCtrl_isSigned <= entriesNext_3_aluCtrl_isSigned;
    entries_3_aluCtrl_logicOp <= entriesNext_3_aluCtrl_logicOp;
    entries_3_shiftCtrl_valid <= entriesNext_3_shiftCtrl_valid;
    entries_3_shiftCtrl_isRight <= entriesNext_3_shiftCtrl_isRight;
    entries_3_shiftCtrl_isArithmetic <= entriesNext_3_shiftCtrl_isArithmetic;
    entries_3_shiftCtrl_isRotate <= entriesNext_3_shiftCtrl_isRotate;
    entries_3_shiftCtrl_isDoubleWord <= entriesNext_3_shiftCtrl_isDoubleWord;
    entries_3_imm <= entriesNext_3_imm;
    entries_3_immUsage <= entriesNext_3_immUsage;
  end


endmodule

module LA32RSimpleDecoder (
  input  wire [31:0]   io_instruction,
  input  wire [31:0]   io_pcIn,
  output wire [31:0]   io_decodedUop_pc,
  output reg           io_decodedUop_isValid,
  output reg  [4:0]    io_decodedUop_uopCode,
  output reg  [3:0]    io_decodedUop_exeUnit,
  output wire [1:0]    io_decodedUop_isa,
  output reg  [4:0]    io_decodedUop_archDest_idx,
  output reg  [1:0]    io_decodedUop_archDest_rtype,
  output reg           io_decodedUop_writeArchDestEn,
  output reg  [4:0]    io_decodedUop_archSrc1_idx,
  output reg  [1:0]    io_decodedUop_archSrc1_rtype,
  output reg           io_decodedUop_useArchSrc1,
  output reg  [4:0]    io_decodedUop_archSrc2_idx,
  output reg  [1:0]    io_decodedUop_archSrc2_rtype,
  output reg           io_decodedUop_useArchSrc2,
  output wire          io_decodedUop_usePcForAddr,
  output reg  [31:0]   io_decodedUop_imm,
  output reg  [2:0]    io_decodedUop_immUsage,
  output reg           io_decodedUop_aluCtrl_valid,
  output reg           io_decodedUop_aluCtrl_isSub,
  output reg           io_decodedUop_aluCtrl_isAdd,
  output reg           io_decodedUop_aluCtrl_isSigned,
  output reg  [1:0]    io_decodedUop_aluCtrl_logicOp,
  output reg           io_decodedUop_shiftCtrl_valid,
  output reg           io_decodedUop_shiftCtrl_isRight,
  output reg           io_decodedUop_shiftCtrl_isArithmetic,
  output wire          io_decodedUop_shiftCtrl_isRotate,
  output wire          io_decodedUop_shiftCtrl_isDoubleWord,
  output reg           io_decodedUop_mulDivCtrl_valid,
  output wire          io_decodedUop_mulDivCtrl_isDiv,
  output reg           io_decodedUop_mulDivCtrl_isSigned,
  output wire          io_decodedUop_mulDivCtrl_isWordOp,
  output reg  [1:0]    io_decodedUop_memCtrl_size,
  output reg           io_decodedUop_memCtrl_isSignedLoad,
  output reg           io_decodedUop_memCtrl_isStore,
  output wire          io_decodedUop_memCtrl_isLoadLinked,
  output wire          io_decodedUop_memCtrl_isStoreCond,
  output wire [4:0]    io_decodedUop_memCtrl_atomicOp,
  output wire          io_decodedUop_memCtrl_isFence,
  output wire [7:0]    io_decodedUop_memCtrl_fenceMode,
  output wire          io_decodedUop_memCtrl_isCacheOp,
  output wire [4:0]    io_decodedUop_memCtrl_cacheOpType,
  output wire          io_decodedUop_memCtrl_isPrefetch,
  output reg  [4:0]    io_decodedUop_branchCtrl_condition,
  output reg           io_decodedUop_branchCtrl_isJump,
  output reg           io_decodedUop_branchCtrl_isLink,
  output reg  [4:0]    io_decodedUop_branchCtrl_linkReg_idx,
  output wire [1:0]    io_decodedUop_branchCtrl_linkReg_rtype,
  output reg           io_decodedUop_branchCtrl_isIndirect,
  output wire [2:0]    io_decodedUop_branchCtrl_laCfIdx,
  output wire [3:0]    io_decodedUop_fpuCtrl_opType,
  output wire [1:0]    io_decodedUop_fpuCtrl_fpSizeSrc1,
  output wire [1:0]    io_decodedUop_fpuCtrl_fpSizeSrc2,
  output wire [1:0]    io_decodedUop_fpuCtrl_fpSizeDest,
  output wire [2:0]    io_decodedUop_fpuCtrl_roundingMode,
  output wire          io_decodedUop_fpuCtrl_isIntegerDest,
  output wire          io_decodedUop_fpuCtrl_isSignedCvt,
  output wire          io_decodedUop_fpuCtrl_fmaNegSrc1,
  output wire [4:0]    io_decodedUop_fpuCtrl_fcmpCond,
  output wire [13:0]   io_decodedUop_csrCtrl_csrAddr,
  output wire          io_decodedUop_csrCtrl_isWrite,
  output wire          io_decodedUop_csrCtrl_isRead,
  output wire          io_decodedUop_csrCtrl_isExchange,
  output wire          io_decodedUop_csrCtrl_useUimmAsSrc,
  output wire [19:0]   io_decodedUop_sysCtrl_sysCode,
  output wire          io_decodedUop_sysCtrl_isExceptionReturn,
  output wire          io_decodedUop_sysCtrl_isTlbOp,
  output wire [3:0]    io_decodedUop_sysCtrl_tlbOpType,
  output reg  [1:0]    io_decodedUop_decodeExceptionCode,
  output reg           io_decodedUop_hasDecodeException,
  output wire          io_decodedUop_isMicrocode,
  output wire [7:0]    io_decodedUop_microcodeEntry,
  output wire          io_decodedUop_isSerializing,
  output reg           io_decodedUop_isBranchOrJump,
  output wire          io_decodedUop_branchPrediction_isTaken,
  output wire [31:0]   io_decodedUop_branchPrediction_target,
  output wire          io_decodedUop_branchPrediction_wasPredicted
);
  localparam BaseUopCode_NOP = 5'd0;
  localparam BaseUopCode_ILLEGAL = 5'd1;
  localparam BaseUopCode_ALU = 5'd2;
  localparam BaseUopCode_SHIFT = 5'd3;
  localparam BaseUopCode_MUL = 5'd4;
  localparam BaseUopCode_DIV = 5'd5;
  localparam BaseUopCode_LOAD = 5'd6;
  localparam BaseUopCode_STORE = 5'd7;
  localparam BaseUopCode_ATOMIC = 5'd8;
  localparam BaseUopCode_MEM_BARRIER = 5'd9;
  localparam BaseUopCode_PREFETCH = 5'd10;
  localparam BaseUopCode_BRANCH = 5'd11;
  localparam BaseUopCode_JUMP_REG = 5'd12;
  localparam BaseUopCode_JUMP_IMM = 5'd13;
  localparam BaseUopCode_SYSTEM_OP = 5'd14;
  localparam BaseUopCode_CSR_ACCESS = 5'd15;
  localparam BaseUopCode_FPU_ALU = 5'd16;
  localparam BaseUopCode_FPU_CVT = 5'd17;
  localparam BaseUopCode_FPU_CMP = 5'd18;
  localparam BaseUopCode_FPU_SEL = 5'd19;
  localparam BaseUopCode_LA_BITMANIP = 5'd20;
  localparam BaseUopCode_LA_CACOP = 5'd21;
  localparam BaseUopCode_LA_TLB = 5'd22;
  localparam BaseUopCode_IDLE = 5'd23;
  localparam ExeUnitType_NONE = 4'd0;
  localparam ExeUnitType_ALU_INT = 4'd1;
  localparam ExeUnitType_MUL_INT = 4'd2;
  localparam ExeUnitType_DIV_INT = 4'd3;
  localparam ExeUnitType_MEM = 4'd4;
  localparam ExeUnitType_BRU = 4'd5;
  localparam ExeUnitType_CSR = 4'd6;
  localparam ExeUnitType_FPU_ADD_MUL_CVT_CMP = 4'd7;
  localparam ExeUnitType_FPU_DIV_SQRT = 4'd8;
  localparam IsaType_UNKNOWN = 2'd0;
  localparam IsaType_DEMO = 2'd1;
  localparam IsaType_RISCV = 2'd2;
  localparam IsaType_LOONGARCH = 2'd3;
  localparam ArchRegType_GPR = 2'd0;
  localparam ArchRegType_FPR = 2'd1;
  localparam ArchRegType_CSR = 2'd2;
  localparam ArchRegType_LA_CF = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;
  localparam BranchCondition_NUL = 5'd0;
  localparam BranchCondition_EQ = 5'd1;
  localparam BranchCondition_NE = 5'd2;
  localparam BranchCondition_LT = 5'd3;
  localparam BranchCondition_GE = 5'd4;
  localparam BranchCondition_LTU = 5'd5;
  localparam BranchCondition_GEU = 5'd6;
  localparam BranchCondition_EQZ = 5'd7;
  localparam BranchCondition_NEZ = 5'd8;
  localparam BranchCondition_LTZ = 5'd9;
  localparam BranchCondition_GEZ = 5'd10;
  localparam BranchCondition_GTZ = 5'd11;
  localparam BranchCondition_LEZ = 5'd12;
  localparam BranchCondition_F_EQ = 5'd13;
  localparam BranchCondition_F_NE = 5'd14;
  localparam BranchCondition_F_LT = 5'd15;
  localparam BranchCondition_F_LE = 5'd16;
  localparam BranchCondition_F_UN = 5'd17;
  localparam BranchCondition_LA_CF_TRUE = 5'd18;
  localparam BranchCondition_LA_CF_FALSE = 5'd19;
  localparam DecodeExCode_INVALID = 2'd0;
  localparam DecodeExCode_FETCH_ERROR = 2'd1;
  localparam DecodeExCode_DECODE_ERROR = 2'd2;
  localparam DecodeExCode_OK = 2'd3;

  wire       [31:0]   _zz_imm_sext_12;
  wire       [11:0]   _zz_imm_sext_12_1;
  wire       [31:0]   _zz_imm_zext_12;
  wire       [11:0]   _zz_imm_zext_12_1;
  wire       [31:0]   _zz_imm_pcadd_u12i;
  wire       [19:0]   _zz_imm_pcadd_u12i_1;
  wire       [31:0]   _zz_imm_branch_16;
  wire       [17:0]   _zz_imm_branch_16_1;
  wire       [15:0]   _zz_imm_branch_16_2;
  wire       [31:0]   _zz_imm_branch_26;
  wire       [27:0]   _zz_imm_branch_26_1;
  wire       [25:0]   _zz_imm_branch_26_2;
  wire       [31:0]   _zz_imm_shift_5;
  wire       [4:0]    _zz_imm_shift_5_1;
  wire       [31:0]   fields_inst;
  wire       [4:0]    r0_idx;
  wire       [4:0]    r1_idx;
  wire       [31:0]   imm_sext_12;
  wire       [31:0]   imm_zext_12;
  wire       [31:0]   imm_lu12i;
  wire       [31:0]   imm_pcadd_u12i;
  wire       [31:0]   imm_branch_16;
  wire       [31:0]   imm_branch_26;
  wire       [31:0]   imm_shift_5;
  wire                is_add_w;
  wire                is_sub_w;
  wire                is_and;
  wire                is_or;
  wire                is_xor;
  wire                is_mul_w;
  wire                is_sll_w;
  wire                is_srl_w;
  wire                is_sra_w;
  wire                is_slli_w;
  wire                is_srli_w;
  wire                is_srai_w;
  wire                is_addi_w;
  wire                is_slti;
  wire                is_andi;
  wire                is_ori;
  wire                is_ld_b;
  wire                is_ld_w;
  wire                is_st_b;
  wire                is_st_w;
  wire                is_lu12i;
  wire                is_pcaddu12i;
  wire                is_jirl;
  wire                is_b;
  wire                is_bl;
  wire                is_beq;
  wire                is_bne;
  wire                is_bltu;
  wire                is_idle;
  wire                is_r_type_alu;
  wire                is_r_type_shift;
  wire                is_r_type;
  wire                is_shift_imm;
  wire                is_i_type;
  wire                is_load;
  wire                is_store;
  wire                is_mem_op;
  wire                is_branch;
  wire                is_jump;
  wire                is_branch_or_jump;
  wire                isValid;
  wire                when_LA32RSimpleDecoder_l174;
  wire                when_LA32RSimpleDecoder_l175;
  wire                when_LA32RSimpleDecoder_l179;
  wire                when_LA32RSimpleDecoder_l185;
  wire                when_LA32RSimpleDecoder_l199;
  wire                when_LA32RSimpleDecoder_l202;
  wire                when_LA32RSimpleDecoder_l206;
  wire                when_LA32RSimpleDecoder_l216;
  wire                when_LA32RSimpleDecoder_l217;
  wire                when_LA32RSimpleDecoder_l220;
  wire                when_LA32RSimpleDecoder_l221;
  wire                when_LA32RSimpleDecoder_l225;
  wire                when_LA32RSimpleDecoder_l229;
  wire                when_LA32RSimpleDecoder_l236;
  wire                when_LA32RSimpleDecoder_l237;
  wire                when_LA32RSimpleDecoder_l239;
  wire                when_LA32RSimpleDecoder_l240;
  wire                when_LA32RSimpleDecoder_l249;
  wire                when_LA32RSimpleDecoder_l250;
  wire                when_LA32RSimpleDecoder_l260;
  wire                when_LA32RSimpleDecoder_l261;
  wire                when_LA32RSimpleDecoder_l266;
  wire                when_LA32RSimpleDecoder_l275;
  `ifndef SYNTHESIS
  reg [87:0] io_decodedUop_uopCode_string;
  reg [151:0] io_decodedUop_exeUnit_string;
  reg [71:0] io_decodedUop_isa_string;
  reg [39:0] io_decodedUop_archDest_rtype_string;
  reg [39:0] io_decodedUop_archSrc1_rtype_string;
  reg [39:0] io_decodedUop_archSrc2_rtype_string;
  reg [103:0] io_decodedUop_immUsage_string;
  reg [39:0] io_decodedUop_aluCtrl_logicOp_string;
  reg [7:0] io_decodedUop_memCtrl_size_string;
  reg [87:0] io_decodedUop_branchCtrl_condition_string;
  reg [39:0] io_decodedUop_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_decodedUop_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_decodedUop_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_decodedUop_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_decodedUop_decodeExceptionCode_string;
  `endif


  assign _zz_imm_sext_12_1 = fields_inst[21 : 10];
  assign _zz_imm_sext_12 = {{20{_zz_imm_sext_12_1[11]}}, _zz_imm_sext_12_1};
  assign _zz_imm_zext_12_1 = fields_inst[21 : 10];
  assign _zz_imm_zext_12 = {20'd0, _zz_imm_zext_12_1};
  assign _zz_imm_pcadd_u12i = ({12'd0,_zz_imm_pcadd_u12i_1} <<< 4'd12);
  assign _zz_imm_pcadd_u12i_1 = fields_inst[24 : 5];
  assign _zz_imm_branch_16_1 = ({2'd0,_zz_imm_branch_16_2} <<< 2'd2);
  assign _zz_imm_branch_16 = {{14{_zz_imm_branch_16_1[17]}}, _zz_imm_branch_16_1};
  assign _zz_imm_branch_16_2 = fields_inst[25 : 10];
  assign _zz_imm_branch_26_1 = ({2'd0,_zz_imm_branch_26_2} <<< 2'd2);
  assign _zz_imm_branch_26 = {{4{_zz_imm_branch_26_1[27]}}, _zz_imm_branch_26_1};
  assign _zz_imm_branch_26_2 = {fields_inst[25 : 16],fields_inst[15 : 0]};
  assign _zz_imm_shift_5_1 = fields_inst[14 : 10];
  assign _zz_imm_shift_5 = {27'd0, _zz_imm_shift_5_1};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_decodedUop_uopCode)
      BaseUopCode_NOP : io_decodedUop_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_decodedUop_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_decodedUop_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_decodedUop_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_decodedUop_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_decodedUop_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_decodedUop_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_decodedUop_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_decodedUop_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_decodedUop_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_decodedUop_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_decodedUop_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_decodedUop_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_decodedUop_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_decodedUop_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_decodedUop_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_decodedUop_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_decodedUop_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_decodedUop_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_decodedUop_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_decodedUop_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_decodedUop_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_decodedUop_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_decodedUop_uopCode_string = "IDLE       ";
      default : io_decodedUop_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_exeUnit)
      ExeUnitType_NONE : io_decodedUop_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_decodedUop_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_decodedUop_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_decodedUop_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_decodedUop_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_decodedUop_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_decodedUop_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_decodedUop_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_decodedUop_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_decodedUop_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_isa)
      IsaType_UNKNOWN : io_decodedUop_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_decodedUop_isa_string = "DEMO     ";
      IsaType_RISCV : io_decodedUop_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_decodedUop_isa_string = "LOONGARCH";
      default : io_decodedUop_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_archDest_rtype)
      ArchRegType_GPR : io_decodedUop_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_decodedUop_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_decodedUop_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_decodedUop_archDest_rtype_string = "LA_CF";
      default : io_decodedUop_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_archSrc1_rtype)
      ArchRegType_GPR : io_decodedUop_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_decodedUop_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_decodedUop_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_decodedUop_archSrc1_rtype_string = "LA_CF";
      default : io_decodedUop_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_archSrc2_rtype)
      ArchRegType_GPR : io_decodedUop_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_decodedUop_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_decodedUop_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_decodedUop_archSrc2_rtype_string = "LA_CF";
      default : io_decodedUop_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_immUsage)
      ImmUsageType_NONE : io_decodedUop_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_decodedUop_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_decodedUop_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_decodedUop_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_decodedUop_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_decodedUop_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_decodedUop_immUsage_string = "JUMP_OFFSET  ";
      default : io_decodedUop_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_aluCtrl_logicOp)
      LogicOp_NONE : io_decodedUop_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_decodedUop_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_decodedUop_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_decodedUop_aluCtrl_logicOp_string = "XOR_1";
      default : io_decodedUop_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_memCtrl_size)
      MemAccessSize_B : io_decodedUop_memCtrl_size_string = "B";
      MemAccessSize_H : io_decodedUop_memCtrl_size_string = "H";
      MemAccessSize_W : io_decodedUop_memCtrl_size_string = "W";
      MemAccessSize_D : io_decodedUop_memCtrl_size_string = "D";
      default : io_decodedUop_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_branchCtrl_condition)
      BranchCondition_NUL : io_decodedUop_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_decodedUop_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_decodedUop_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_decodedUop_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_decodedUop_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_decodedUop_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_decodedUop_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_decodedUop_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_decodedUop_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_decodedUop_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_decodedUop_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_decodedUop_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_decodedUop_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_decodedUop_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_decodedUop_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_decodedUop_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_decodedUop_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_decodedUop_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_decodedUop_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_decodedUop_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_decodedUop_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_decodedUop_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_decodedUop_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_decodedUop_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_decodedUop_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_decodedUop_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_decodedUop_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_decodedUop_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_decodedUop_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_decodedUop_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_decodedUop_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_decodedUop_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_decodedUop_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_decodedUop_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_decodedUop_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_decodedUop_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_decodedUop_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_decodedUop_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_decodedUop_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_decodedUop_fpuCtrl_fpSizeDest_string = "D";
      default : io_decodedUop_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_decodedUop_decodeExceptionCode)
      DecodeExCode_INVALID : io_decodedUop_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_decodedUop_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_decodedUop_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_decodedUop_decodeExceptionCode_string = "OK          ";
      default : io_decodedUop_decodeExceptionCode_string = "????????????";
    endcase
  end
  `endif

  assign fields_inst = io_instruction;
  assign r0_idx = 5'h0;
  assign r1_idx = 5'h01;
  assign imm_sext_12 = _zz_imm_sext_12;
  assign imm_zext_12 = _zz_imm_zext_12;
  assign imm_lu12i = {fields_inst[24 : 5],12'h0};
  assign imm_pcadd_u12i = _zz_imm_pcadd_u12i;
  assign imm_branch_16 = _zz_imm_branch_16;
  assign imm_branch_26 = _zz_imm_branch_26;
  assign imm_shift_5 = _zz_imm_shift_5;
  assign is_add_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h020));
  assign is_sub_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h022));
  assign is_and = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h029));
  assign is_or = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h02a));
  assign is_xor = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h02b));
  assign is_mul_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h038));
  assign is_sll_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h02e));
  assign is_srl_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h02f));
  assign is_sra_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h030));
  assign is_slli_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h081));
  assign is_srli_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h089));
  assign is_srai_w = ((fields_inst[31 : 25] == 7'h0) && (fields_inst[24 : 15] == 10'h091));
  assign is_addi_w = ((fields_inst[31 : 25] == 7'h01) && (fields_inst[24 : 22] == 3'b010));
  assign is_slti = ((fields_inst[31 : 25] == 7'h01) && (fields_inst[24 : 22] == 3'b000));
  assign is_andi = ((fields_inst[31 : 25] == 7'h01) && (fields_inst[24 : 22] == 3'b101));
  assign is_ori = ((fields_inst[31 : 25] == 7'h01) && (fields_inst[24 : 22] == 3'b110));
  assign is_ld_b = ((fields_inst[31 : 25] == 7'h14) && (fields_inst[24 : 22] == 3'b000));
  assign is_ld_w = ((fields_inst[31 : 25] == 7'h14) && (fields_inst[24 : 22] == 3'b010));
  assign is_st_b = ((fields_inst[31 : 25] == 7'h14) && (fields_inst[24 : 22] == 3'b100));
  assign is_st_w = ((fields_inst[31 : 25] == 7'h14) && (fields_inst[24 : 22] == 3'b110));
  assign is_lu12i = (fields_inst[31 : 25] == 7'h0a);
  assign is_pcaddu12i = (fields_inst[31 : 25] == 7'h0e);
  assign is_jirl = (fields_inst[31 : 26] == 6'h13);
  assign is_b = (fields_inst[31 : 26] == 6'h14);
  assign is_bl = (fields_inst[31 : 26] == 6'h15);
  assign is_beq = (fields_inst[31 : 26] == 6'h16);
  assign is_bne = (fields_inst[31 : 26] == 6'h17);
  assign is_bltu = (fields_inst[31 : 26] == 6'h1a);
  assign is_idle = ((fields_inst[31 : 25] == 7'h03) && (fields_inst[24 : 15] == 10'h091));
  assign is_r_type_alu = ((((is_add_w || is_sub_w) || is_and) || is_or) || is_xor);
  assign is_r_type_shift = ((is_sll_w || is_srl_w) || is_sra_w);
  assign is_r_type = ((is_r_type_alu || is_r_type_shift) || is_mul_w);
  assign is_shift_imm = ((is_slli_w || is_srli_w) || is_srai_w);
  assign is_i_type = (((is_addi_w || is_slti) || is_andi) || is_ori);
  assign is_load = (is_ld_b || is_ld_w);
  assign is_store = (is_st_b || is_st_w);
  assign is_mem_op = (is_load || is_store);
  assign is_branch = ((is_beq || is_bne) || is_bltu);
  assign is_jump = ((is_b || is_bl) || is_jirl);
  assign is_branch_or_jump = (is_branch || is_jump);
  assign io_decodedUop_pc = io_pcIn;
  always @(*) begin
    io_decodedUop_isValid = 1'b0;
    io_decodedUop_isValid = isValid;
  end

  always @(*) begin
    io_decodedUop_uopCode = BaseUopCode_NOP;
    io_decodedUop_uopCode = BaseUopCode_ILLEGAL;
    if(when_LA32RSimpleDecoder_l174) begin
      io_decodedUop_uopCode = BaseUopCode_ALU;
    end
    if(when_LA32RSimpleDecoder_l175) begin
      io_decodedUop_uopCode = BaseUopCode_SHIFT;
    end
    if(is_mul_w) begin
      io_decodedUop_uopCode = BaseUopCode_MUL;
    end
    if(is_load) begin
      io_decodedUop_uopCode = BaseUopCode_LOAD;
    end
    if(is_store) begin
      io_decodedUop_uopCode = BaseUopCode_STORE;
    end
    if(when_LA32RSimpleDecoder_l179) begin
      io_decodedUop_uopCode = BaseUopCode_JUMP_IMM;
    end
    if(is_jirl) begin
      io_decodedUop_uopCode = BaseUopCode_JUMP_REG;
    end
    if(is_branch) begin
      io_decodedUop_uopCode = BaseUopCode_BRANCH;
    end
    if(is_idle) begin
      io_decodedUop_uopCode = BaseUopCode_IDLE;
    end
    if(when_LA32RSimpleDecoder_l275) begin
      io_decodedUop_uopCode = BaseUopCode_ILLEGAL;
    end
  end

  always @(*) begin
    io_decodedUop_exeUnit = ExeUnitType_NONE;
    io_decodedUop_exeUnit = ExeUnitType_NONE;
    if(when_LA32RSimpleDecoder_l185) begin
      io_decodedUop_exeUnit = ExeUnitType_ALU_INT;
    end
    if(is_mul_w) begin
      io_decodedUop_exeUnit = ExeUnitType_MUL_INT;
    end
    if(is_mem_op) begin
      io_decodedUop_exeUnit = ExeUnitType_MEM;
    end
    if(is_branch_or_jump) begin
      io_decodedUop_exeUnit = ExeUnitType_BRU;
    end
  end

  assign io_decodedUop_isa = IsaType_LOONGARCH;
  always @(*) begin
    io_decodedUop_archDest_idx = 5'h0;
    io_decodedUop_archDest_idx = 5'h0;
    if(when_LA32RSimpleDecoder_l202) begin
      io_decodedUop_archDest_idx = fields_inst[4 : 0];
    end
    if(is_bl) begin
      io_decodedUop_archDest_idx = r1_idx;
    end
  end

  always @(*) begin
    io_decodedUop_archDest_rtype = ArchRegType_GPR;
    if(io_decodedUop_writeArchDestEn) begin
      io_decodedUop_archDest_rtype = ArchRegType_GPR;
    end
  end

  always @(*) begin
    io_decodedUop_writeArchDestEn = 1'b0;
    io_decodedUop_writeArchDestEn = 1'b0;
    if(when_LA32RSimpleDecoder_l206) begin
      io_decodedUop_writeArchDestEn = 1'b1;
    end
    if(is_bl) begin
      io_decodedUop_writeArchDestEn = 1'b1;
    end
  end

  always @(*) begin
    io_decodedUop_archSrc1_idx = 5'h0;
    io_decodedUop_archSrc1_idx = 5'h0;
    if(io_decodedUop_useArchSrc1) begin
      io_decodedUop_archSrc1_idx = fields_inst[9 : 5];
    end
  end

  always @(*) begin
    io_decodedUop_archSrc1_rtype = ArchRegType_GPR;
    if(io_decodedUop_useArchSrc1) begin
      io_decodedUop_archSrc1_rtype = ArchRegType_GPR;
    end
  end

  always @(*) begin
    io_decodedUop_useArchSrc1 = 1'b0;
    io_decodedUop_useArchSrc1 = (((((is_r_type || is_shift_imm) || is_i_type) || is_mem_op) || is_jirl) || is_branch);
  end

  always @(*) begin
    io_decodedUop_archSrc2_idx = 5'h0;
    io_decodedUop_archSrc2_idx = 5'h0;
    if(is_r_type) begin
      io_decodedUop_archSrc2_idx = fields_inst[14 : 10];
    end
    if(when_LA32RSimpleDecoder_l199) begin
      io_decodedUop_archSrc2_idx = fields_inst[4 : 0];
    end
  end

  always @(*) begin
    io_decodedUop_archSrc2_rtype = ArchRegType_GPR;
    if(io_decodedUop_useArchSrc2) begin
      io_decodedUop_archSrc2_rtype = ArchRegType_GPR;
    end
  end

  always @(*) begin
    io_decodedUop_useArchSrc2 = 1'b0;
    io_decodedUop_useArchSrc2 = ((is_r_type || is_store) || is_branch);
  end

  assign io_decodedUop_usePcForAddr = 1'b0;
  always @(*) begin
    io_decodedUop_imm = 32'h0;
    io_decodedUop_imm = 32'h0;
    if(when_LA32RSimpleDecoder_l216) begin
      io_decodedUop_imm = imm_sext_12;
    end
    if(when_LA32RSimpleDecoder_l217) begin
      io_decodedUop_imm = imm_zext_12;
    end
    if(is_lu12i) begin
      io_decodedUop_imm = imm_lu12i;
    end
    if(is_pcaddu12i) begin
      io_decodedUop_imm = imm_pcadd_u12i;
    end
    if(when_LA32RSimpleDecoder_l220) begin
      io_decodedUop_imm = imm_branch_16;
    end
    if(when_LA32RSimpleDecoder_l221) begin
      io_decodedUop_imm = imm_branch_26;
    end
    if(is_shift_imm) begin
      io_decodedUop_imm = imm_shift_5;
    end
  end

  always @(*) begin
    io_decodedUop_immUsage = ImmUsageType_NONE;
    io_decodedUop_immUsage = ImmUsageType_NONE;
    if(when_LA32RSimpleDecoder_l225) begin
      io_decodedUop_immUsage = ImmUsageType_SRC_ALU;
    end
    if(is_shift_imm) begin
      io_decodedUop_immUsage = ImmUsageType_SRC_SHIFT_AMT;
    end
    if(is_mem_op) begin
      io_decodedUop_immUsage = ImmUsageType_MEM_OFFSET;
    end
    if(is_branch) begin
      io_decodedUop_immUsage = ImmUsageType_BRANCH_OFFSET;
    end
    if(when_LA32RSimpleDecoder_l229) begin
      io_decodedUop_immUsage = ImmUsageType_JUMP_OFFSET;
    end
    if(is_jirl) begin
      io_decodedUop_immUsage = ImmUsageType_BRANCH_OFFSET;
    end
  end

  always @(*) begin
    io_decodedUop_aluCtrl_valid = 1'b0;
    io_decodedUop_aluCtrl_valid = (((((((is_add_w || is_addi_w) || is_lu12i) || is_pcaddu12i) || (is_sub_w || is_slti)) || (is_and || is_andi)) || (is_or || is_ori)) || is_xor);
  end

  always @(*) begin
    io_decodedUop_aluCtrl_isSub = 1'b0;
    if(when_LA32RSimpleDecoder_l237) begin
      io_decodedUop_aluCtrl_isSub = 1'b1;
    end
  end

  always @(*) begin
    io_decodedUop_aluCtrl_isAdd = 1'b0;
    if(when_LA32RSimpleDecoder_l236) begin
      io_decodedUop_aluCtrl_isAdd = 1'b1;
    end
  end

  always @(*) begin
    io_decodedUop_aluCtrl_isSigned = 1'b0;
    if(is_slti) begin
      io_decodedUop_aluCtrl_isSigned = 1'b1;
    end
  end

  always @(*) begin
    io_decodedUop_aluCtrl_logicOp = LogicOp_NONE;
    if(when_LA32RSimpleDecoder_l239) begin
      io_decodedUop_aluCtrl_logicOp = LogicOp_AND_1;
    end
    if(when_LA32RSimpleDecoder_l240) begin
      io_decodedUop_aluCtrl_logicOp = LogicOp_OR_1;
    end
    if(is_xor) begin
      io_decodedUop_aluCtrl_logicOp = LogicOp_XOR_1;
    end
  end

  always @(*) begin
    io_decodedUop_shiftCtrl_valid = 1'b0;
    io_decodedUop_shiftCtrl_valid = (((is_srl_w || is_srli_w) || is_sra_w) || is_srai_w);
  end

  always @(*) begin
    io_decodedUop_shiftCtrl_isRight = 1'b0;
    if(when_LA32RSimpleDecoder_l249) begin
      io_decodedUop_shiftCtrl_isRight = 1'b1;
    end
  end

  always @(*) begin
    io_decodedUop_shiftCtrl_isArithmetic = 1'b0;
    if(when_LA32RSimpleDecoder_l250) begin
      io_decodedUop_shiftCtrl_isArithmetic = 1'b1;
    end
  end

  assign io_decodedUop_shiftCtrl_isRotate = 1'b0;
  assign io_decodedUop_shiftCtrl_isDoubleWord = 1'b0;
  always @(*) begin
    io_decodedUop_mulDivCtrl_valid = 1'b0;
    io_decodedUop_mulDivCtrl_valid = is_mul_w;
  end

  assign io_decodedUop_mulDivCtrl_isDiv = 1'b0;
  always @(*) begin
    io_decodedUop_mulDivCtrl_isSigned = 1'b0;
    if(is_mul_w) begin
      io_decodedUop_mulDivCtrl_isSigned = 1'b1;
    end
  end

  assign io_decodedUop_mulDivCtrl_isWordOp = 1'b0;
  always @(*) begin
    io_decodedUop_memCtrl_size = MemAccessSize_W;
    if(when_LA32RSimpleDecoder_l260) begin
      io_decodedUop_memCtrl_size = MemAccessSize_B;
    end
    if(when_LA32RSimpleDecoder_l261) begin
      io_decodedUop_memCtrl_size = MemAccessSize_W;
    end
  end

  always @(*) begin
    io_decodedUop_memCtrl_isSignedLoad = 1'b0;
    if(is_load) begin
      io_decodedUop_memCtrl_isSignedLoad = 1'b1;
    end
  end

  always @(*) begin
    io_decodedUop_memCtrl_isStore = 1'b0;
    if(is_store) begin
      io_decodedUop_memCtrl_isStore = 1'b1;
    end
  end

  assign io_decodedUop_memCtrl_isLoadLinked = 1'b0;
  assign io_decodedUop_memCtrl_isStoreCond = 1'b0;
  assign io_decodedUop_memCtrl_atomicOp = 5'h0;
  assign io_decodedUop_memCtrl_isFence = 1'b0;
  assign io_decodedUop_memCtrl_fenceMode = 8'h0;
  assign io_decodedUop_memCtrl_isCacheOp = 1'b0;
  assign io_decodedUop_memCtrl_cacheOpType = 5'h0;
  assign io_decodedUop_memCtrl_isPrefetch = 1'b0;
  always @(*) begin
    io_decodedUop_branchCtrl_condition = BranchCondition_NUL;
    if(is_beq) begin
      io_decodedUop_branchCtrl_condition = BranchCondition_EQ;
    end
    if(is_bne) begin
      io_decodedUop_branchCtrl_condition = BranchCondition_NE;
    end
    if(is_bltu) begin
      io_decodedUop_branchCtrl_condition = BranchCondition_LTU;
    end
  end

  always @(*) begin
    io_decodedUop_branchCtrl_isJump = 1'b0;
    if(is_jump) begin
      io_decodedUop_branchCtrl_isJump = 1'b1;
    end
  end

  always @(*) begin
    io_decodedUop_branchCtrl_isLink = 1'b0;
    if(when_LA32RSimpleDecoder_l266) begin
      io_decodedUop_branchCtrl_isLink = 1'b1;
    end
  end

  always @(*) begin
    io_decodedUop_branchCtrl_linkReg_idx = 5'h0;
    if(is_bl) begin
      io_decodedUop_branchCtrl_linkReg_idx = r1_idx;
    end
    if(is_jirl) begin
      io_decodedUop_branchCtrl_linkReg_idx = fields_inst[4 : 0];
    end
  end

  assign io_decodedUop_branchCtrl_linkReg_rtype = ArchRegType_GPR;
  always @(*) begin
    io_decodedUop_branchCtrl_isIndirect = 1'b0;
    if(is_jirl) begin
      io_decodedUop_branchCtrl_isIndirect = 1'b1;
    end
  end

  assign io_decodedUop_branchCtrl_laCfIdx = 3'b000;
  assign io_decodedUop_fpuCtrl_opType = 4'b0000;
  assign io_decodedUop_fpuCtrl_fpSizeSrc1 = MemAccessSize_W;
  assign io_decodedUop_fpuCtrl_fpSizeSrc2 = MemAccessSize_W;
  assign io_decodedUop_fpuCtrl_fpSizeDest = MemAccessSize_W;
  assign io_decodedUop_fpuCtrl_roundingMode = 3'b000;
  assign io_decodedUop_fpuCtrl_isIntegerDest = 1'b0;
  assign io_decodedUop_fpuCtrl_isSignedCvt = 1'b0;
  assign io_decodedUop_fpuCtrl_fmaNegSrc1 = 1'b0;
  assign io_decodedUop_fpuCtrl_fcmpCond = 5'h0;
  assign io_decodedUop_csrCtrl_csrAddr = 14'h0;
  assign io_decodedUop_csrCtrl_isWrite = 1'b0;
  assign io_decodedUop_csrCtrl_isRead = 1'b0;
  assign io_decodedUop_csrCtrl_isExchange = 1'b0;
  assign io_decodedUop_csrCtrl_useUimmAsSrc = 1'b0;
  assign io_decodedUop_sysCtrl_sysCode = 20'h0;
  assign io_decodedUop_sysCtrl_isExceptionReturn = 1'b0;
  assign io_decodedUop_sysCtrl_isTlbOp = 1'b0;
  assign io_decodedUop_sysCtrl_tlbOpType = 4'b0000;
  always @(*) begin
    io_decodedUop_decodeExceptionCode = DecodeExCode_OK;
    if(when_LA32RSimpleDecoder_l275) begin
      io_decodedUop_decodeExceptionCode = DecodeExCode_DECODE_ERROR;
    end
  end

  always @(*) begin
    io_decodedUop_hasDecodeException = 1'b0;
    if(when_LA32RSimpleDecoder_l275) begin
      io_decodedUop_hasDecodeException = 1'b1;
    end
  end

  assign io_decodedUop_isMicrocode = 1'b0;
  assign io_decodedUop_microcodeEntry = 8'h0;
  assign io_decodedUop_isSerializing = 1'b0;
  always @(*) begin
    io_decodedUop_isBranchOrJump = 1'b0;
    io_decodedUop_isBranchOrJump = is_branch_or_jump;
  end

  assign io_decodedUop_branchPrediction_isTaken = 1'b0;
  assign io_decodedUop_branchPrediction_target = 32'h0;
  assign io_decodedUop_branchPrediction_wasPredicted = 1'b0;
  assign isValid = (((((((is_r_type || is_shift_imm) || is_i_type) || is_mem_op) || is_lu12i) || is_pcaddu12i) || is_branch_or_jump) || is_idle);
  assign when_LA32RSimpleDecoder_l174 = (((is_r_type_alu || is_i_type) || is_lu12i) || is_pcaddu12i);
  assign when_LA32RSimpleDecoder_l175 = (is_r_type_shift || is_shift_imm);
  assign when_LA32RSimpleDecoder_l179 = (is_b || is_bl);
  assign when_LA32RSimpleDecoder_l185 = (((((is_r_type || is_shift_imm) || is_i_type) || is_lu12i) || is_pcaddu12i) || is_idle);
  assign when_LA32RSimpleDecoder_l199 = (is_store || is_branch);
  assign when_LA32RSimpleDecoder_l202 = ((((((is_r_type || is_shift_imm) || is_i_type) || is_load) || is_lu12i) || is_pcaddu12i) || is_jirl);
  assign when_LA32RSimpleDecoder_l206 = (((((((is_r_type || is_shift_imm) || is_i_type) || is_load) || is_lu12i) || is_pcaddu12i) || is_jirl) && (fields_inst[4 : 0] != r0_idx));
  assign when_LA32RSimpleDecoder_l216 = ((is_addi_w || is_slti) || is_mem_op);
  assign when_LA32RSimpleDecoder_l217 = (is_andi || is_ori);
  assign when_LA32RSimpleDecoder_l220 = (is_branch || is_jirl);
  assign when_LA32RSimpleDecoder_l221 = (is_b || is_bl);
  assign when_LA32RSimpleDecoder_l225 = ((is_i_type || is_lu12i) || is_pcaddu12i);
  assign when_LA32RSimpleDecoder_l229 = (is_b || is_bl);
  assign when_LA32RSimpleDecoder_l236 = (((is_add_w || is_addi_w) || is_lu12i) || is_pcaddu12i);
  assign when_LA32RSimpleDecoder_l237 = (is_sub_w || is_slti);
  assign when_LA32RSimpleDecoder_l239 = (is_and || is_andi);
  assign when_LA32RSimpleDecoder_l240 = (is_or || is_ori);
  assign when_LA32RSimpleDecoder_l249 = (((is_srl_w || is_srli_w) || is_sra_w) || is_srai_w);
  assign when_LA32RSimpleDecoder_l250 = (is_sra_w || is_srai_w);
  assign when_LA32RSimpleDecoder_l260 = (is_ld_b || is_st_b);
  assign when_LA32RSimpleDecoder_l261 = (is_ld_w || is_st_w);
  assign when_LA32RSimpleDecoder_l266 = (is_bl || is_jirl);
  assign when_LA32RSimpleDecoder_l275 = (! isValid);

endmodule

//OneShot_6 replaced by OneShot

//OneShot_5 replaced by OneShot

module StreamArbiter_6 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [5:0]    io_inputs_0_payload_physRegIdx,
  input  wire [31:0]   io_inputs_0_payload_physRegData,
  input  wire [3:0]    io_inputs_0_payload_robPtr,
  input  wire          io_inputs_0_payload_isFPR,
  input  wire          io_inputs_0_payload_hasException,
  input  wire [7:0]    io_inputs_0_payload_exceptionCode,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [5:0]    io_inputs_1_payload_physRegIdx,
  input  wire [31:0]   io_inputs_1_payload_physRegData,
  input  wire [3:0]    io_inputs_1_payload_robPtr,
  input  wire          io_inputs_1_payload_isFPR,
  input  wire          io_inputs_1_payload_hasException,
  input  wire [7:0]    io_inputs_1_payload_exceptionCode,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [5:0]    io_inputs_2_payload_physRegIdx,
  input  wire [31:0]   io_inputs_2_payload_physRegData,
  input  wire [3:0]    io_inputs_2_payload_robPtr,
  input  wire          io_inputs_2_payload_isFPR,
  input  wire          io_inputs_2_payload_hasException,
  input  wire [7:0]    io_inputs_2_payload_exceptionCode,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [5:0]    io_output_payload_physRegIdx,
  output wire [31:0]   io_output_payload_physRegData,
  output wire [3:0]    io_output_payload_robPtr,
  output wire          io_output_payload_isFPR,
  output wire          io_output_payload_hasException,
  output wire [7:0]    io_output_payload_exceptionCode,
  output wire [1:0]    io_chosen,
  output wire [2:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [5:0]    _zz__zz_maskProposal_0_2;
  wire       [5:0]    _zz__zz_maskProposal_0_2_1;
  wire       [2:0]    _zz__zz_maskProposal_0_2_2;
  reg        [5:0]    _zz_io_output_payload_physRegIdx_1;
  reg        [31:0]   _zz_io_output_payload_physRegData;
  reg        [3:0]    _zz_io_output_payload_robPtr;
  reg                 _zz_io_output_payload_isFPR;
  reg                 _zz_io_output_payload_hasException;
  reg        [7:0]    _zz_io_output_payload_exceptionCode;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire       [2:0]    _zz_maskProposal_0;
  wire       [5:0]    _zz_maskProposal_0_1;
  wire       [5:0]    _zz_maskProposal_0_2;
  wire       [2:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire       [1:0]    _zz_io_output_payload_physRegIdx;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_1,{maskLocked_0,maskLocked_2}};
  assign _zz__zz_maskProposal_0_2_1 = {3'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(_zz_io_output_payload_physRegIdx)
      2'b00 : begin
        _zz_io_output_payload_physRegIdx_1 = io_inputs_0_payload_physRegIdx;
        _zz_io_output_payload_physRegData = io_inputs_0_payload_physRegData;
        _zz_io_output_payload_robPtr = io_inputs_0_payload_robPtr;
        _zz_io_output_payload_isFPR = io_inputs_0_payload_isFPR;
        _zz_io_output_payload_hasException = io_inputs_0_payload_hasException;
        _zz_io_output_payload_exceptionCode = io_inputs_0_payload_exceptionCode;
      end
      2'b01 : begin
        _zz_io_output_payload_physRegIdx_1 = io_inputs_1_payload_physRegIdx;
        _zz_io_output_payload_physRegData = io_inputs_1_payload_physRegData;
        _zz_io_output_payload_robPtr = io_inputs_1_payload_robPtr;
        _zz_io_output_payload_isFPR = io_inputs_1_payload_isFPR;
        _zz_io_output_payload_hasException = io_inputs_1_payload_hasException;
        _zz_io_output_payload_exceptionCode = io_inputs_1_payload_exceptionCode;
      end
      default : begin
        _zz_io_output_payload_physRegIdx_1 = io_inputs_2_payload_physRegIdx;
        _zz_io_output_payload_physRegData = io_inputs_2_payload_physRegData;
        _zz_io_output_payload_robPtr = io_inputs_2_payload_robPtr;
        _zz_io_output_payload_isFPR = io_inputs_2_payload_isFPR;
        _zz_io_output_payload_hasException = io_inputs_2_payload_hasException;
        _zz_io_output_payload_exceptionCode = io_inputs_2_payload_exceptionCode;
      end
    endcase
  end

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign _zz_maskProposal_0 = {io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[5 : 3] | _zz_maskProposal_0_2[2 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2));
  assign _zz_io_output_payload_physRegIdx = {maskRouted_2,maskRouted_1};
  assign io_output_payload_physRegIdx = _zz_io_output_payload_physRegIdx_1;
  assign io_output_payload_physRegData = _zz_io_output_payload_physRegData;
  assign io_output_payload_robPtr = _zz_io_output_payload_robPtr;
  assign io_output_payload_isFPR = _zz_io_output_payload_isFPR;
  assign io_output_payload_hasException = _zz_io_output_payload_hasException;
  assign io_output_payload_exceptionCode = _zz_io_output_payload_exceptionCode;
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_inputs_1_ready = ((1'b0 || maskRouted_1) && io_output_ready);
  assign io_inputs_2_ready = ((1'b0 || maskRouted_2) && io_output_ready);
  assign io_chosenOH = {maskRouted_2,{maskRouted_1,maskRouted_0}};
  assign _zz_io_chosen = io_chosenOH[1];
  assign _zz_io_chosen_1 = io_chosenOH[2];
  assign io_chosen = {_zz_io_chosen_1,_zz_io_chosen};
  always @(posedge clk) begin
    if(reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module EightSegmentDisplayController (
  input  wire [7:0]    io_value,
  input  wire          io_dp0,
  input  wire          io_dp1,
  output wire [7:0]    io_dpy0_out,
  output wire [7:0]    io_dpy1_out
);

  wire       [3:0]    displayArea_digit0;
  wire       [3:0]    displayArea_digit1;
  reg        [6:0]    displayArea_seg0;
  reg        [6:0]    displayArea_seg1;

  assign displayArea_digit0 = io_value[3 : 0];
  assign displayArea_digit1 = io_value[7 : 4];
  always @(*) begin
    case(displayArea_digit0)
      4'b0000 : begin
        displayArea_seg0 = 7'h3f;
      end
      4'b0001 : begin
        displayArea_seg0 = 7'h09;
      end
      4'b0010 : begin
        displayArea_seg0 = 7'h5e;
      end
      4'b0011 : begin
        displayArea_seg0 = 7'h5b;
      end
      4'b0100 : begin
        displayArea_seg0 = 7'h69;
      end
      4'b0101 : begin
        displayArea_seg0 = 7'h73;
      end
      4'b0110 : begin
        displayArea_seg0 = 7'h77;
      end
      4'b0111 : begin
        displayArea_seg0 = 7'h19;
      end
      4'b1000 : begin
        displayArea_seg0 = 7'h7f;
      end
      4'b1001 : begin
        displayArea_seg0 = 7'h7b;
      end
      4'b1010 : begin
        displayArea_seg0 = 7'h7d;
      end
      4'b1011 : begin
        displayArea_seg0 = 7'h67;
      end
      4'b1100 : begin
        displayArea_seg0 = 7'h36;
      end
      4'b1101 : begin
        displayArea_seg0 = 7'h4f;
      end
      4'b1110 : begin
        displayArea_seg0 = 7'h76;
      end
      default : begin
        displayArea_seg0 = 7'h74;
      end
    endcase
  end

  always @(*) begin
    case(displayArea_digit1)
      4'b0000 : begin
        displayArea_seg1 = 7'h3f;
      end
      4'b0001 : begin
        displayArea_seg1 = 7'h09;
      end
      4'b0010 : begin
        displayArea_seg1 = 7'h5e;
      end
      4'b0011 : begin
        displayArea_seg1 = 7'h5b;
      end
      4'b0100 : begin
        displayArea_seg1 = 7'h69;
      end
      4'b0101 : begin
        displayArea_seg1 = 7'h73;
      end
      4'b0110 : begin
        displayArea_seg1 = 7'h77;
      end
      4'b0111 : begin
        displayArea_seg1 = 7'h19;
      end
      4'b1000 : begin
        displayArea_seg1 = 7'h7f;
      end
      4'b1001 : begin
        displayArea_seg1 = 7'h7b;
      end
      4'b1010 : begin
        displayArea_seg1 = 7'h7d;
      end
      4'b1011 : begin
        displayArea_seg1 = 7'h67;
      end
      4'b1100 : begin
        displayArea_seg1 = 7'h36;
      end
      4'b1101 : begin
        displayArea_seg1 = 7'h4f;
      end
      4'b1110 : begin
        displayArea_seg1 = 7'h76;
      end
      default : begin
        displayArea_seg1 = 7'h74;
      end
    endcase
  end

  assign io_dpy0_out = {displayArea_seg0,io_dp0};
  assign io_dpy1_out = {displayArea_seg1,io_dp1};

endmodule

module RenameUnit (
  input  wire [31:0]   io_decodedUopsIn_0_pc,
  input  wire          io_decodedUopsIn_0_isValid,
  input  wire [4:0]    io_decodedUopsIn_0_uopCode,
  input  wire [3:0]    io_decodedUopsIn_0_exeUnit,
  input  wire [1:0]    io_decodedUopsIn_0_isa,
  input  wire [4:0]    io_decodedUopsIn_0_archDest_idx,
  input  wire [1:0]    io_decodedUopsIn_0_archDest_rtype,
  input  wire          io_decodedUopsIn_0_writeArchDestEn,
  input  wire [4:0]    io_decodedUopsIn_0_archSrc1_idx,
  input  wire [1:0]    io_decodedUopsIn_0_archSrc1_rtype,
  input  wire          io_decodedUopsIn_0_useArchSrc1,
  input  wire [4:0]    io_decodedUopsIn_0_archSrc2_idx,
  input  wire [1:0]    io_decodedUopsIn_0_archSrc2_rtype,
  input  wire          io_decodedUopsIn_0_useArchSrc2,
  input  wire          io_decodedUopsIn_0_usePcForAddr,
  input  wire [31:0]   io_decodedUopsIn_0_imm,
  input  wire [2:0]    io_decodedUopsIn_0_immUsage,
  input  wire          io_decodedUopsIn_0_aluCtrl_valid,
  input  wire          io_decodedUopsIn_0_aluCtrl_isSub,
  input  wire          io_decodedUopsIn_0_aluCtrl_isAdd,
  input  wire          io_decodedUopsIn_0_aluCtrl_isSigned,
  input  wire [1:0]    io_decodedUopsIn_0_aluCtrl_logicOp,
  input  wire          io_decodedUopsIn_0_shiftCtrl_valid,
  input  wire          io_decodedUopsIn_0_shiftCtrl_isRight,
  input  wire          io_decodedUopsIn_0_shiftCtrl_isArithmetic,
  input  wire          io_decodedUopsIn_0_shiftCtrl_isRotate,
  input  wire          io_decodedUopsIn_0_shiftCtrl_isDoubleWord,
  input  wire          io_decodedUopsIn_0_mulDivCtrl_valid,
  input  wire          io_decodedUopsIn_0_mulDivCtrl_isDiv,
  input  wire          io_decodedUopsIn_0_mulDivCtrl_isSigned,
  input  wire          io_decodedUopsIn_0_mulDivCtrl_isWordOp,
  input  wire [1:0]    io_decodedUopsIn_0_memCtrl_size,
  input  wire          io_decodedUopsIn_0_memCtrl_isSignedLoad,
  input  wire          io_decodedUopsIn_0_memCtrl_isStore,
  input  wire          io_decodedUopsIn_0_memCtrl_isLoadLinked,
  input  wire          io_decodedUopsIn_0_memCtrl_isStoreCond,
  input  wire [4:0]    io_decodedUopsIn_0_memCtrl_atomicOp,
  input  wire          io_decodedUopsIn_0_memCtrl_isFence,
  input  wire [7:0]    io_decodedUopsIn_0_memCtrl_fenceMode,
  input  wire          io_decodedUopsIn_0_memCtrl_isCacheOp,
  input  wire [4:0]    io_decodedUopsIn_0_memCtrl_cacheOpType,
  input  wire          io_decodedUopsIn_0_memCtrl_isPrefetch,
  input  wire [4:0]    io_decodedUopsIn_0_branchCtrl_condition,
  input  wire          io_decodedUopsIn_0_branchCtrl_isJump,
  input  wire          io_decodedUopsIn_0_branchCtrl_isLink,
  input  wire [4:0]    io_decodedUopsIn_0_branchCtrl_linkReg_idx,
  input  wire [1:0]    io_decodedUopsIn_0_branchCtrl_linkReg_rtype,
  input  wire          io_decodedUopsIn_0_branchCtrl_isIndirect,
  input  wire [2:0]    io_decodedUopsIn_0_branchCtrl_laCfIdx,
  input  wire [3:0]    io_decodedUopsIn_0_fpuCtrl_opType,
  input  wire [1:0]    io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1,
  input  wire [1:0]    io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2,
  input  wire [1:0]    io_decodedUopsIn_0_fpuCtrl_fpSizeDest,
  input  wire [2:0]    io_decodedUopsIn_0_fpuCtrl_roundingMode,
  input  wire          io_decodedUopsIn_0_fpuCtrl_isIntegerDest,
  input  wire          io_decodedUopsIn_0_fpuCtrl_isSignedCvt,
  input  wire          io_decodedUopsIn_0_fpuCtrl_fmaNegSrc1,
  input  wire [4:0]    io_decodedUopsIn_0_fpuCtrl_fcmpCond,
  input  wire [13:0]   io_decodedUopsIn_0_csrCtrl_csrAddr,
  input  wire          io_decodedUopsIn_0_csrCtrl_isWrite,
  input  wire          io_decodedUopsIn_0_csrCtrl_isRead,
  input  wire          io_decodedUopsIn_0_csrCtrl_isExchange,
  input  wire          io_decodedUopsIn_0_csrCtrl_useUimmAsSrc,
  input  wire [19:0]   io_decodedUopsIn_0_sysCtrl_sysCode,
  input  wire          io_decodedUopsIn_0_sysCtrl_isExceptionReturn,
  input  wire          io_decodedUopsIn_0_sysCtrl_isTlbOp,
  input  wire [3:0]    io_decodedUopsIn_0_sysCtrl_tlbOpType,
  input  wire [1:0]    io_decodedUopsIn_0_decodeExceptionCode,
  input  wire          io_decodedUopsIn_0_hasDecodeException,
  input  wire          io_decodedUopsIn_0_isMicrocode,
  input  wire [7:0]    io_decodedUopsIn_0_microcodeEntry,
  input  wire          io_decodedUopsIn_0_isSerializing,
  input  wire          io_decodedUopsIn_0_isBranchOrJump,
  input  wire          io_decodedUopsIn_0_branchPrediction_isTaken,
  input  wire [31:0]   io_decodedUopsIn_0_branchPrediction_target,
  input  wire          io_decodedUopsIn_0_branchPrediction_wasPredicted,
  input  wire [5:0]    io_physRegsIn_0,
  output wire [31:0]   io_renamedUopsOut_0_decoded_pc,
  output wire          io_renamedUopsOut_0_decoded_isValid,
  output wire [4:0]    io_renamedUopsOut_0_decoded_uopCode,
  output wire [3:0]    io_renamedUopsOut_0_decoded_exeUnit,
  output wire [1:0]    io_renamedUopsOut_0_decoded_isa,
  output wire [4:0]    io_renamedUopsOut_0_decoded_archDest_idx,
  output wire [1:0]    io_renamedUopsOut_0_decoded_archDest_rtype,
  output wire          io_renamedUopsOut_0_decoded_writeArchDestEn,
  output wire [4:0]    io_renamedUopsOut_0_decoded_archSrc1_idx,
  output wire [1:0]    io_renamedUopsOut_0_decoded_archSrc1_rtype,
  output wire          io_renamedUopsOut_0_decoded_useArchSrc1,
  output wire [4:0]    io_renamedUopsOut_0_decoded_archSrc2_idx,
  output wire [1:0]    io_renamedUopsOut_0_decoded_archSrc2_rtype,
  output wire          io_renamedUopsOut_0_decoded_useArchSrc2,
  output wire          io_renamedUopsOut_0_decoded_usePcForAddr,
  output wire [31:0]   io_renamedUopsOut_0_decoded_imm,
  output wire [2:0]    io_renamedUopsOut_0_decoded_immUsage,
  output wire          io_renamedUopsOut_0_decoded_aluCtrl_valid,
  output wire          io_renamedUopsOut_0_decoded_aluCtrl_isSub,
  output wire          io_renamedUopsOut_0_decoded_aluCtrl_isAdd,
  output wire          io_renamedUopsOut_0_decoded_aluCtrl_isSigned,
  output wire [1:0]    io_renamedUopsOut_0_decoded_aluCtrl_logicOp,
  output wire          io_renamedUopsOut_0_decoded_shiftCtrl_valid,
  output wire          io_renamedUopsOut_0_decoded_shiftCtrl_isRight,
  output wire          io_renamedUopsOut_0_decoded_shiftCtrl_isArithmetic,
  output wire          io_renamedUopsOut_0_decoded_shiftCtrl_isRotate,
  output wire          io_renamedUopsOut_0_decoded_shiftCtrl_isDoubleWord,
  output wire          io_renamedUopsOut_0_decoded_mulDivCtrl_valid,
  output wire          io_renamedUopsOut_0_decoded_mulDivCtrl_isDiv,
  output wire          io_renamedUopsOut_0_decoded_mulDivCtrl_isSigned,
  output wire          io_renamedUopsOut_0_decoded_mulDivCtrl_isWordOp,
  output wire [1:0]    io_renamedUopsOut_0_decoded_memCtrl_size,
  output wire          io_renamedUopsOut_0_decoded_memCtrl_isSignedLoad,
  output wire          io_renamedUopsOut_0_decoded_memCtrl_isStore,
  output wire          io_renamedUopsOut_0_decoded_memCtrl_isLoadLinked,
  output wire          io_renamedUopsOut_0_decoded_memCtrl_isStoreCond,
  output wire [4:0]    io_renamedUopsOut_0_decoded_memCtrl_atomicOp,
  output wire          io_renamedUopsOut_0_decoded_memCtrl_isFence,
  output wire [7:0]    io_renamedUopsOut_0_decoded_memCtrl_fenceMode,
  output wire          io_renamedUopsOut_0_decoded_memCtrl_isCacheOp,
  output wire [4:0]    io_renamedUopsOut_0_decoded_memCtrl_cacheOpType,
  output wire          io_renamedUopsOut_0_decoded_memCtrl_isPrefetch,
  output wire [4:0]    io_renamedUopsOut_0_decoded_branchCtrl_condition,
  output wire          io_renamedUopsOut_0_decoded_branchCtrl_isJump,
  output wire          io_renamedUopsOut_0_decoded_branchCtrl_isLink,
  output wire [4:0]    io_renamedUopsOut_0_decoded_branchCtrl_linkReg_idx,
  output wire [1:0]    io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype,
  output wire          io_renamedUopsOut_0_decoded_branchCtrl_isIndirect,
  output wire [2:0]    io_renamedUopsOut_0_decoded_branchCtrl_laCfIdx,
  output wire [3:0]    io_renamedUopsOut_0_decoded_fpuCtrl_opType,
  output wire [1:0]    io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1,
  output wire [1:0]    io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2,
  output wire [1:0]    io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest,
  output wire [2:0]    io_renamedUopsOut_0_decoded_fpuCtrl_roundingMode,
  output wire          io_renamedUopsOut_0_decoded_fpuCtrl_isIntegerDest,
  output wire          io_renamedUopsOut_0_decoded_fpuCtrl_isSignedCvt,
  output wire          io_renamedUopsOut_0_decoded_fpuCtrl_fmaNegSrc1,
  output wire [4:0]    io_renamedUopsOut_0_decoded_fpuCtrl_fcmpCond,
  output wire [13:0]   io_renamedUopsOut_0_decoded_csrCtrl_csrAddr,
  output wire          io_renamedUopsOut_0_decoded_csrCtrl_isWrite,
  output wire          io_renamedUopsOut_0_decoded_csrCtrl_isRead,
  output wire          io_renamedUopsOut_0_decoded_csrCtrl_isExchange,
  output wire          io_renamedUopsOut_0_decoded_csrCtrl_useUimmAsSrc,
  output wire [19:0]   io_renamedUopsOut_0_decoded_sysCtrl_sysCode,
  output wire          io_renamedUopsOut_0_decoded_sysCtrl_isExceptionReturn,
  output wire          io_renamedUopsOut_0_decoded_sysCtrl_isTlbOp,
  output wire [3:0]    io_renamedUopsOut_0_decoded_sysCtrl_tlbOpType,
  output wire [1:0]    io_renamedUopsOut_0_decoded_decodeExceptionCode,
  output wire          io_renamedUopsOut_0_decoded_hasDecodeException,
  output wire          io_renamedUopsOut_0_decoded_isMicrocode,
  output wire [7:0]    io_renamedUopsOut_0_decoded_microcodeEntry,
  output wire          io_renamedUopsOut_0_decoded_isSerializing,
  output wire          io_renamedUopsOut_0_decoded_isBranchOrJump,
  output wire          io_renamedUopsOut_0_decoded_branchPrediction_isTaken,
  output wire [31:0]   io_renamedUopsOut_0_decoded_branchPrediction_target,
  output wire          io_renamedUopsOut_0_decoded_branchPrediction_wasPredicted,
  output wire [5:0]    io_renamedUopsOut_0_rename_physSrc1_idx,
  output wire          io_renamedUopsOut_0_rename_physSrc1IsFpr,
  output wire [5:0]    io_renamedUopsOut_0_rename_physSrc2_idx,
  output wire          io_renamedUopsOut_0_rename_physSrc2IsFpr,
  output reg  [5:0]    io_renamedUopsOut_0_rename_physDest_idx,
  output reg           io_renamedUopsOut_0_rename_physDestIsFpr,
  output reg  [5:0]    io_renamedUopsOut_0_rename_oldPhysDest_idx,
  output reg           io_renamedUopsOut_0_rename_oldPhysDestIsFpr,
  output reg           io_renamedUopsOut_0_rename_allocatesPhysDest,
  output reg           io_renamedUopsOut_0_rename_writesToPhysReg,
  output wire [3:0]    io_renamedUopsOut_0_robPtr,
  output wire [15:0]   io_renamedUopsOut_0_uniqueId,
  output wire          io_renamedUopsOut_0_dispatched,
  output wire          io_renamedUopsOut_0_executed,
  output wire          io_renamedUopsOut_0_hasException,
  output wire [7:0]    io_renamedUopsOut_0_exceptionCode,
  output wire [0:0]    io_numPhysRegsRequired,
  output wire [4:0]    io_ratReadPorts_0_archReg,
  input  wire [5:0]    io_ratReadPorts_0_physReg,
  output wire [4:0]    io_ratReadPorts_1_archReg,
  input  wire [5:0]    io_ratReadPorts_1_physReg,
  output wire [4:0]    io_ratReadPorts_2_archReg,
  input  wire [5:0]    io_ratReadPorts_2_physReg,
  output wire          io_ratWritePorts_0_wen,
  output wire [4:0]    io_ratWritePorts_0_archReg,
  output wire [5:0]    io_ratWritePorts_0_physReg,
  input  wire          clk,
  input  wire          reset
);
  localparam BaseUopCode_NOP = 5'd0;
  localparam BaseUopCode_ILLEGAL = 5'd1;
  localparam BaseUopCode_ALU = 5'd2;
  localparam BaseUopCode_SHIFT = 5'd3;
  localparam BaseUopCode_MUL = 5'd4;
  localparam BaseUopCode_DIV = 5'd5;
  localparam BaseUopCode_LOAD = 5'd6;
  localparam BaseUopCode_STORE = 5'd7;
  localparam BaseUopCode_ATOMIC = 5'd8;
  localparam BaseUopCode_MEM_BARRIER = 5'd9;
  localparam BaseUopCode_PREFETCH = 5'd10;
  localparam BaseUopCode_BRANCH = 5'd11;
  localparam BaseUopCode_JUMP_REG = 5'd12;
  localparam BaseUopCode_JUMP_IMM = 5'd13;
  localparam BaseUopCode_SYSTEM_OP = 5'd14;
  localparam BaseUopCode_CSR_ACCESS = 5'd15;
  localparam BaseUopCode_FPU_ALU = 5'd16;
  localparam BaseUopCode_FPU_CVT = 5'd17;
  localparam BaseUopCode_FPU_CMP = 5'd18;
  localparam BaseUopCode_FPU_SEL = 5'd19;
  localparam BaseUopCode_LA_BITMANIP = 5'd20;
  localparam BaseUopCode_LA_CACOP = 5'd21;
  localparam BaseUopCode_LA_TLB = 5'd22;
  localparam BaseUopCode_IDLE = 5'd23;
  localparam ExeUnitType_NONE = 4'd0;
  localparam ExeUnitType_ALU_INT = 4'd1;
  localparam ExeUnitType_MUL_INT = 4'd2;
  localparam ExeUnitType_DIV_INT = 4'd3;
  localparam ExeUnitType_MEM = 4'd4;
  localparam ExeUnitType_BRU = 4'd5;
  localparam ExeUnitType_CSR = 4'd6;
  localparam ExeUnitType_FPU_ADD_MUL_CVT_CMP = 4'd7;
  localparam ExeUnitType_FPU_DIV_SQRT = 4'd8;
  localparam IsaType_UNKNOWN = 2'd0;
  localparam IsaType_DEMO = 2'd1;
  localparam IsaType_RISCV = 2'd2;
  localparam IsaType_LOONGARCH = 2'd3;
  localparam ArchRegType_GPR = 2'd0;
  localparam ArchRegType_FPR = 2'd1;
  localparam ArchRegType_CSR = 2'd2;
  localparam ArchRegType_LA_CF = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;
  localparam BranchCondition_NUL = 5'd0;
  localparam BranchCondition_EQ = 5'd1;
  localparam BranchCondition_NE = 5'd2;
  localparam BranchCondition_LT = 5'd3;
  localparam BranchCondition_GE = 5'd4;
  localparam BranchCondition_LTU = 5'd5;
  localparam BranchCondition_GEU = 5'd6;
  localparam BranchCondition_EQZ = 5'd7;
  localparam BranchCondition_NEZ = 5'd8;
  localparam BranchCondition_LTZ = 5'd9;
  localparam BranchCondition_GEZ = 5'd10;
  localparam BranchCondition_GTZ = 5'd11;
  localparam BranchCondition_LEZ = 5'd12;
  localparam BranchCondition_F_EQ = 5'd13;
  localparam BranchCondition_F_NE = 5'd14;
  localparam BranchCondition_F_LT = 5'd15;
  localparam BranchCondition_F_LE = 5'd16;
  localparam BranchCondition_F_UN = 5'd17;
  localparam BranchCondition_LA_CF_TRUE = 5'd18;
  localparam BranchCondition_LA_CF_FALSE = 5'd19;
  localparam DecodeExCode_INVALID = 2'd0;
  localparam DecodeExCode_FETCH_ERROR = 2'd1;
  localparam DecodeExCode_DECODE_ERROR = 2'd2;
  localparam DecodeExCode_OK = 2'd3;

  wire                uopNeedsNewPhysDest;
  wire                _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [4:0]    toplevel_RenamePlugin_setup_renameUnit_debugDecodedArchSrc2;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg                 toplevel_RenamePlugin_setup_renameUnit_debugDecodedUseArchSrc2;
  (* MARK_DEBUG = "TRUE" , DONT_TOUCH = "TRUE" *) reg        [5:0]    toplevel_RenamePlugin_setup_renameUnit_debugRenamedPhysSrc2;
  `ifndef SYNTHESIS
  reg [87:0] io_decodedUopsIn_0_uopCode_string;
  reg [151:0] io_decodedUopsIn_0_exeUnit_string;
  reg [71:0] io_decodedUopsIn_0_isa_string;
  reg [39:0] io_decodedUopsIn_0_archDest_rtype_string;
  reg [39:0] io_decodedUopsIn_0_archSrc1_rtype_string;
  reg [39:0] io_decodedUopsIn_0_archSrc2_rtype_string;
  reg [103:0] io_decodedUopsIn_0_immUsage_string;
  reg [39:0] io_decodedUopsIn_0_aluCtrl_logicOp_string;
  reg [7:0] io_decodedUopsIn_0_memCtrl_size_string;
  reg [87:0] io_decodedUopsIn_0_branchCtrl_condition_string;
  reg [39:0] io_decodedUopsIn_0_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_decodedUopsIn_0_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_decodedUopsIn_0_decodeExceptionCode_string;
  reg [87:0] io_renamedUopsOut_0_decoded_uopCode_string;
  reg [151:0] io_renamedUopsOut_0_decoded_exeUnit_string;
  reg [71:0] io_renamedUopsOut_0_decoded_isa_string;
  reg [39:0] io_renamedUopsOut_0_decoded_archDest_rtype_string;
  reg [39:0] io_renamedUopsOut_0_decoded_archSrc1_rtype_string;
  reg [39:0] io_renamedUopsOut_0_decoded_archSrc2_rtype_string;
  reg [103:0] io_renamedUopsOut_0_decoded_immUsage_string;
  reg [39:0] io_renamedUopsOut_0_decoded_aluCtrl_logicOp_string;
  reg [7:0] io_renamedUopsOut_0_decoded_memCtrl_size_string;
  reg [87:0] io_renamedUopsOut_0_decoded_branchCtrl_condition_string;
  reg [39:0] io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_renamedUopsOut_0_decoded_decodeExceptionCode_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_decodedUopsIn_0_uopCode)
      BaseUopCode_NOP : io_decodedUopsIn_0_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_decodedUopsIn_0_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_decodedUopsIn_0_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_decodedUopsIn_0_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_decodedUopsIn_0_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_decodedUopsIn_0_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_decodedUopsIn_0_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_decodedUopsIn_0_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_decodedUopsIn_0_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_decodedUopsIn_0_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_decodedUopsIn_0_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_decodedUopsIn_0_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_decodedUopsIn_0_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_decodedUopsIn_0_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_decodedUopsIn_0_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_decodedUopsIn_0_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_decodedUopsIn_0_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_decodedUopsIn_0_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_decodedUopsIn_0_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_decodedUopsIn_0_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_decodedUopsIn_0_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_decodedUopsIn_0_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_decodedUopsIn_0_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_decodedUopsIn_0_uopCode_string = "IDLE       ";
      default : io_decodedUopsIn_0_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_exeUnit)
      ExeUnitType_NONE : io_decodedUopsIn_0_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_decodedUopsIn_0_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_decodedUopsIn_0_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_decodedUopsIn_0_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_decodedUopsIn_0_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_decodedUopsIn_0_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_decodedUopsIn_0_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_decodedUopsIn_0_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_decodedUopsIn_0_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_decodedUopsIn_0_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_isa)
      IsaType_UNKNOWN : io_decodedUopsIn_0_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_decodedUopsIn_0_isa_string = "DEMO     ";
      IsaType_RISCV : io_decodedUopsIn_0_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_decodedUopsIn_0_isa_string = "LOONGARCH";
      default : io_decodedUopsIn_0_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_archDest_rtype)
      ArchRegType_GPR : io_decodedUopsIn_0_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_decodedUopsIn_0_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_decodedUopsIn_0_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_decodedUopsIn_0_archDest_rtype_string = "LA_CF";
      default : io_decodedUopsIn_0_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_archSrc1_rtype)
      ArchRegType_GPR : io_decodedUopsIn_0_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_decodedUopsIn_0_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_decodedUopsIn_0_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_decodedUopsIn_0_archSrc1_rtype_string = "LA_CF";
      default : io_decodedUopsIn_0_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_archSrc2_rtype)
      ArchRegType_GPR : io_decodedUopsIn_0_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_decodedUopsIn_0_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_decodedUopsIn_0_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_decodedUopsIn_0_archSrc2_rtype_string = "LA_CF";
      default : io_decodedUopsIn_0_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_immUsage)
      ImmUsageType_NONE : io_decodedUopsIn_0_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_decodedUopsIn_0_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_decodedUopsIn_0_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_decodedUopsIn_0_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_decodedUopsIn_0_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_decodedUopsIn_0_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_decodedUopsIn_0_immUsage_string = "JUMP_OFFSET  ";
      default : io_decodedUopsIn_0_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_aluCtrl_logicOp)
      LogicOp_NONE : io_decodedUopsIn_0_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_decodedUopsIn_0_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_decodedUopsIn_0_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_decodedUopsIn_0_aluCtrl_logicOp_string = "XOR_1";
      default : io_decodedUopsIn_0_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_memCtrl_size)
      MemAccessSize_B : io_decodedUopsIn_0_memCtrl_size_string = "B";
      MemAccessSize_H : io_decodedUopsIn_0_memCtrl_size_string = "H";
      MemAccessSize_W : io_decodedUopsIn_0_memCtrl_size_string = "W";
      MemAccessSize_D : io_decodedUopsIn_0_memCtrl_size_string = "D";
      default : io_decodedUopsIn_0_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_branchCtrl_condition)
      BranchCondition_NUL : io_decodedUopsIn_0_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_decodedUopsIn_0_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_decodedUopsIn_0_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_decodedUopsIn_0_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_decodedUopsIn_0_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_decodedUopsIn_0_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_decodedUopsIn_0_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_decodedUopsIn_0_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_decodedUopsIn_0_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_decodedUopsIn_0_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_decodedUopsIn_0_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_decodedUopsIn_0_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_decodedUopsIn_0_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_decodedUopsIn_0_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_decodedUopsIn_0_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_decodedUopsIn_0_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_decodedUopsIn_0_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_decodedUopsIn_0_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_decodedUopsIn_0_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_decodedUopsIn_0_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_decodedUopsIn_0_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_decodedUopsIn_0_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_decodedUopsIn_0_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_decodedUopsIn_0_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_decodedUopsIn_0_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_decodedUopsIn_0_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_decodedUopsIn_0_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_decodedUopsIn_0_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_decodedUopsIn_0_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_decodedUopsIn_0_fpuCtrl_fpSizeDest_string = "D";
      default : io_decodedUopsIn_0_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_decodedUopsIn_0_decodeExceptionCode)
      DecodeExCode_INVALID : io_decodedUopsIn_0_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_decodedUopsIn_0_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_decodedUopsIn_0_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_decodedUopsIn_0_decodeExceptionCode_string = "OK          ";
      default : io_decodedUopsIn_0_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_uopCode)
      BaseUopCode_NOP : io_renamedUopsOut_0_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_renamedUopsOut_0_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_renamedUopsOut_0_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_renamedUopsOut_0_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_renamedUopsOut_0_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_renamedUopsOut_0_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_renamedUopsOut_0_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_renamedUopsOut_0_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_renamedUopsOut_0_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_renamedUopsOut_0_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_renamedUopsOut_0_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_renamedUopsOut_0_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_renamedUopsOut_0_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_renamedUopsOut_0_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_renamedUopsOut_0_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_renamedUopsOut_0_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_renamedUopsOut_0_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_renamedUopsOut_0_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_renamedUopsOut_0_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_renamedUopsOut_0_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_renamedUopsOut_0_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_renamedUopsOut_0_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_renamedUopsOut_0_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_renamedUopsOut_0_decoded_uopCode_string = "IDLE       ";
      default : io_renamedUopsOut_0_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_exeUnit)
      ExeUnitType_NONE : io_renamedUopsOut_0_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_renamedUopsOut_0_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_renamedUopsOut_0_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_renamedUopsOut_0_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_renamedUopsOut_0_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_renamedUopsOut_0_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_renamedUopsOut_0_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_renamedUopsOut_0_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_renamedUopsOut_0_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_renamedUopsOut_0_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_isa)
      IsaType_UNKNOWN : io_renamedUopsOut_0_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_renamedUopsOut_0_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : io_renamedUopsOut_0_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_renamedUopsOut_0_decoded_isa_string = "LOONGARCH";
      default : io_renamedUopsOut_0_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_archDest_rtype)
      ArchRegType_GPR : io_renamedUopsOut_0_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_renamedUopsOut_0_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_renamedUopsOut_0_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_renamedUopsOut_0_decoded_archDest_rtype_string = "LA_CF";
      default : io_renamedUopsOut_0_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_archSrc1_rtype)
      ArchRegType_GPR : io_renamedUopsOut_0_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_renamedUopsOut_0_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_renamedUopsOut_0_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_renamedUopsOut_0_decoded_archSrc1_rtype_string = "LA_CF";
      default : io_renamedUopsOut_0_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_archSrc2_rtype)
      ArchRegType_GPR : io_renamedUopsOut_0_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_renamedUopsOut_0_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_renamedUopsOut_0_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_renamedUopsOut_0_decoded_archSrc2_rtype_string = "LA_CF";
      default : io_renamedUopsOut_0_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_immUsage)
      ImmUsageType_NONE : io_renamedUopsOut_0_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_renamedUopsOut_0_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_renamedUopsOut_0_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_renamedUopsOut_0_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_renamedUopsOut_0_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_renamedUopsOut_0_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_renamedUopsOut_0_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : io_renamedUopsOut_0_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_aluCtrl_logicOp)
      LogicOp_NONE : io_renamedUopsOut_0_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_renamedUopsOut_0_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_renamedUopsOut_0_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_renamedUopsOut_0_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : io_renamedUopsOut_0_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_memCtrl_size)
      MemAccessSize_B : io_renamedUopsOut_0_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : io_renamedUopsOut_0_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : io_renamedUopsOut_0_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : io_renamedUopsOut_0_decoded_memCtrl_size_string = "D";
      default : io_renamedUopsOut_0_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_branchCtrl_condition)
      BranchCondition_NUL : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_renamedUopsOut_0_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_renamedUopsOut_0_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : io_renamedUopsOut_0_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_renamedUopsOut_0_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_renamedUopsOut_0_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_renamedUopsOut_0_decoded_decodeExceptionCode_string = "OK          ";
      default : io_renamedUopsOut_0_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  `endif

  assign uopNeedsNewPhysDest = ((io_decodedUopsIn_0_isValid && io_decodedUopsIn_0_writeArchDestEn) && ((io_decodedUopsIn_0_archDest_rtype == ArchRegType_GPR) || (io_decodedUopsIn_0_archDest_rtype == ArchRegType_FPR)));
  assign io_numPhysRegsRequired = uopNeedsNewPhysDest;
  assign io_ratReadPorts_0_archReg = (io_decodedUopsIn_0_useArchSrc1 ? io_decodedUopsIn_0_archSrc1_idx : 5'h0);
  assign io_ratReadPorts_1_archReg = (io_decodedUopsIn_0_useArchSrc2 ? io_decodedUopsIn_0_archSrc2_idx : 5'h0);
  assign io_ratReadPorts_2_archReg = (uopNeedsNewPhysDest ? io_decodedUopsIn_0_archDest_idx : 5'h0);
  assign io_renamedUopsOut_0_decoded_pc = io_decodedUopsIn_0_pc;
  assign io_renamedUopsOut_0_decoded_isValid = io_decodedUopsIn_0_isValid;
  assign io_renamedUopsOut_0_decoded_uopCode = io_decodedUopsIn_0_uopCode;
  assign io_renamedUopsOut_0_decoded_exeUnit = io_decodedUopsIn_0_exeUnit;
  assign io_renamedUopsOut_0_decoded_isa = io_decodedUopsIn_0_isa;
  assign io_renamedUopsOut_0_decoded_archDest_idx = io_decodedUopsIn_0_archDest_idx;
  assign io_renamedUopsOut_0_decoded_archDest_rtype = io_decodedUopsIn_0_archDest_rtype;
  assign io_renamedUopsOut_0_decoded_writeArchDestEn = io_decodedUopsIn_0_writeArchDestEn;
  assign io_renamedUopsOut_0_decoded_archSrc1_idx = io_decodedUopsIn_0_archSrc1_idx;
  assign io_renamedUopsOut_0_decoded_archSrc1_rtype = io_decodedUopsIn_0_archSrc1_rtype;
  assign io_renamedUopsOut_0_decoded_useArchSrc1 = io_decodedUopsIn_0_useArchSrc1;
  assign io_renamedUopsOut_0_decoded_archSrc2_idx = io_decodedUopsIn_0_archSrc2_idx;
  assign io_renamedUopsOut_0_decoded_archSrc2_rtype = io_decodedUopsIn_0_archSrc2_rtype;
  assign io_renamedUopsOut_0_decoded_useArchSrc2 = io_decodedUopsIn_0_useArchSrc2;
  assign io_renamedUopsOut_0_decoded_usePcForAddr = io_decodedUopsIn_0_usePcForAddr;
  assign io_renamedUopsOut_0_decoded_imm = io_decodedUopsIn_0_imm;
  assign io_renamedUopsOut_0_decoded_immUsage = io_decodedUopsIn_0_immUsage;
  assign io_renamedUopsOut_0_decoded_aluCtrl_valid = io_decodedUopsIn_0_aluCtrl_valid;
  assign io_renamedUopsOut_0_decoded_aluCtrl_isSub = io_decodedUopsIn_0_aluCtrl_isSub;
  assign io_renamedUopsOut_0_decoded_aluCtrl_isAdd = io_decodedUopsIn_0_aluCtrl_isAdd;
  assign io_renamedUopsOut_0_decoded_aluCtrl_isSigned = io_decodedUopsIn_0_aluCtrl_isSigned;
  assign io_renamedUopsOut_0_decoded_aluCtrl_logicOp = io_decodedUopsIn_0_aluCtrl_logicOp;
  assign io_renamedUopsOut_0_decoded_shiftCtrl_valid = io_decodedUopsIn_0_shiftCtrl_valid;
  assign io_renamedUopsOut_0_decoded_shiftCtrl_isRight = io_decodedUopsIn_0_shiftCtrl_isRight;
  assign io_renamedUopsOut_0_decoded_shiftCtrl_isArithmetic = io_decodedUopsIn_0_shiftCtrl_isArithmetic;
  assign io_renamedUopsOut_0_decoded_shiftCtrl_isRotate = io_decodedUopsIn_0_shiftCtrl_isRotate;
  assign io_renamedUopsOut_0_decoded_shiftCtrl_isDoubleWord = io_decodedUopsIn_0_shiftCtrl_isDoubleWord;
  assign io_renamedUopsOut_0_decoded_mulDivCtrl_valid = io_decodedUopsIn_0_mulDivCtrl_valid;
  assign io_renamedUopsOut_0_decoded_mulDivCtrl_isDiv = io_decodedUopsIn_0_mulDivCtrl_isDiv;
  assign io_renamedUopsOut_0_decoded_mulDivCtrl_isSigned = io_decodedUopsIn_0_mulDivCtrl_isSigned;
  assign io_renamedUopsOut_0_decoded_mulDivCtrl_isWordOp = io_decodedUopsIn_0_mulDivCtrl_isWordOp;
  assign io_renamedUopsOut_0_decoded_memCtrl_size = io_decodedUopsIn_0_memCtrl_size;
  assign io_renamedUopsOut_0_decoded_memCtrl_isSignedLoad = io_decodedUopsIn_0_memCtrl_isSignedLoad;
  assign io_renamedUopsOut_0_decoded_memCtrl_isStore = io_decodedUopsIn_0_memCtrl_isStore;
  assign io_renamedUopsOut_0_decoded_memCtrl_isLoadLinked = io_decodedUopsIn_0_memCtrl_isLoadLinked;
  assign io_renamedUopsOut_0_decoded_memCtrl_isStoreCond = io_decodedUopsIn_0_memCtrl_isStoreCond;
  assign io_renamedUopsOut_0_decoded_memCtrl_atomicOp = io_decodedUopsIn_0_memCtrl_atomicOp;
  assign io_renamedUopsOut_0_decoded_memCtrl_isFence = io_decodedUopsIn_0_memCtrl_isFence;
  assign io_renamedUopsOut_0_decoded_memCtrl_fenceMode = io_decodedUopsIn_0_memCtrl_fenceMode;
  assign io_renamedUopsOut_0_decoded_memCtrl_isCacheOp = io_decodedUopsIn_0_memCtrl_isCacheOp;
  assign io_renamedUopsOut_0_decoded_memCtrl_cacheOpType = io_decodedUopsIn_0_memCtrl_cacheOpType;
  assign io_renamedUopsOut_0_decoded_memCtrl_isPrefetch = io_decodedUopsIn_0_memCtrl_isPrefetch;
  assign io_renamedUopsOut_0_decoded_branchCtrl_condition = io_decodedUopsIn_0_branchCtrl_condition;
  assign io_renamedUopsOut_0_decoded_branchCtrl_isJump = io_decodedUopsIn_0_branchCtrl_isJump;
  assign io_renamedUopsOut_0_decoded_branchCtrl_isLink = io_decodedUopsIn_0_branchCtrl_isLink;
  assign io_renamedUopsOut_0_decoded_branchCtrl_linkReg_idx = io_decodedUopsIn_0_branchCtrl_linkReg_idx;
  assign io_renamedUopsOut_0_decoded_branchCtrl_linkReg_rtype = io_decodedUopsIn_0_branchCtrl_linkReg_rtype;
  assign io_renamedUopsOut_0_decoded_branchCtrl_isIndirect = io_decodedUopsIn_0_branchCtrl_isIndirect;
  assign io_renamedUopsOut_0_decoded_branchCtrl_laCfIdx = io_decodedUopsIn_0_branchCtrl_laCfIdx;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_opType = io_decodedUopsIn_0_fpuCtrl_opType;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc1 = io_decodedUopsIn_0_fpuCtrl_fpSizeSrc1;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeSrc2 = io_decodedUopsIn_0_fpuCtrl_fpSizeSrc2;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_fpSizeDest = io_decodedUopsIn_0_fpuCtrl_fpSizeDest;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_roundingMode = io_decodedUopsIn_0_fpuCtrl_roundingMode;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_isIntegerDest = io_decodedUopsIn_0_fpuCtrl_isIntegerDest;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_isSignedCvt = io_decodedUopsIn_0_fpuCtrl_isSignedCvt;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_fmaNegSrc1 = io_decodedUopsIn_0_fpuCtrl_fmaNegSrc1;
  assign io_renamedUopsOut_0_decoded_fpuCtrl_fcmpCond = io_decodedUopsIn_0_fpuCtrl_fcmpCond;
  assign io_renamedUopsOut_0_decoded_csrCtrl_csrAddr = io_decodedUopsIn_0_csrCtrl_csrAddr;
  assign io_renamedUopsOut_0_decoded_csrCtrl_isWrite = io_decodedUopsIn_0_csrCtrl_isWrite;
  assign io_renamedUopsOut_0_decoded_csrCtrl_isRead = io_decodedUopsIn_0_csrCtrl_isRead;
  assign io_renamedUopsOut_0_decoded_csrCtrl_isExchange = io_decodedUopsIn_0_csrCtrl_isExchange;
  assign io_renamedUopsOut_0_decoded_csrCtrl_useUimmAsSrc = io_decodedUopsIn_0_csrCtrl_useUimmAsSrc;
  assign io_renamedUopsOut_0_decoded_sysCtrl_sysCode = io_decodedUopsIn_0_sysCtrl_sysCode;
  assign io_renamedUopsOut_0_decoded_sysCtrl_isExceptionReturn = io_decodedUopsIn_0_sysCtrl_isExceptionReturn;
  assign io_renamedUopsOut_0_decoded_sysCtrl_isTlbOp = io_decodedUopsIn_0_sysCtrl_isTlbOp;
  assign io_renamedUopsOut_0_decoded_sysCtrl_tlbOpType = io_decodedUopsIn_0_sysCtrl_tlbOpType;
  assign io_renamedUopsOut_0_decoded_decodeExceptionCode = io_decodedUopsIn_0_decodeExceptionCode;
  assign io_renamedUopsOut_0_decoded_hasDecodeException = io_decodedUopsIn_0_hasDecodeException;
  assign io_renamedUopsOut_0_decoded_isMicrocode = io_decodedUopsIn_0_isMicrocode;
  assign io_renamedUopsOut_0_decoded_microcodeEntry = io_decodedUopsIn_0_microcodeEntry;
  assign io_renamedUopsOut_0_decoded_isSerializing = io_decodedUopsIn_0_isSerializing;
  assign io_renamedUopsOut_0_decoded_isBranchOrJump = io_decodedUopsIn_0_isBranchOrJump;
  assign io_renamedUopsOut_0_decoded_branchPrediction_isTaken = io_decodedUopsIn_0_branchPrediction_isTaken;
  assign io_renamedUopsOut_0_decoded_branchPrediction_target = io_decodedUopsIn_0_branchPrediction_target;
  assign io_renamedUopsOut_0_decoded_branchPrediction_wasPredicted = io_decodedUopsIn_0_branchPrediction_wasPredicted;
  assign io_renamedUopsOut_0_uniqueId = 16'bxxxxxxxxxxxxxxxx;
  assign io_renamedUopsOut_0_robPtr = 4'bxxxx;
  assign io_renamedUopsOut_0_dispatched = 1'b0;
  assign io_renamedUopsOut_0_executed = 1'b0;
  assign io_renamedUopsOut_0_hasException = 1'b0;
  assign io_renamedUopsOut_0_exceptionCode = 8'h0;
  assign io_renamedUopsOut_0_rename_physSrc1_idx = io_ratReadPorts_0_physReg;
  assign io_renamedUopsOut_0_rename_physSrc1IsFpr = (io_decodedUopsIn_0_archSrc1_rtype == ArchRegType_FPR);
  assign io_renamedUopsOut_0_rename_physSrc2_idx = io_ratReadPorts_1_physReg;
  assign io_renamedUopsOut_0_rename_physSrc2IsFpr = (io_decodedUopsIn_0_archSrc2_rtype == ArchRegType_FPR);
  always @(*) begin
    if(uopNeedsNewPhysDest) begin
      io_renamedUopsOut_0_rename_writesToPhysReg = 1'b1;
    end else begin
      io_renamedUopsOut_0_rename_writesToPhysReg = 1'b0;
    end
  end

  always @(*) begin
    if(uopNeedsNewPhysDest) begin
      io_renamedUopsOut_0_rename_oldPhysDest_idx = io_ratReadPorts_2_physReg;
    end else begin
      io_renamedUopsOut_0_rename_oldPhysDest_idx = 6'h0;
    end
  end

  always @(*) begin
    if(uopNeedsNewPhysDest) begin
      io_renamedUopsOut_0_rename_oldPhysDestIsFpr = (io_decodedUopsIn_0_archDest_rtype == ArchRegType_FPR);
    end else begin
      io_renamedUopsOut_0_rename_oldPhysDestIsFpr = 1'b0;
    end
  end

  always @(*) begin
    if(uopNeedsNewPhysDest) begin
      io_renamedUopsOut_0_rename_allocatesPhysDest = 1'b1;
    end else begin
      io_renamedUopsOut_0_rename_allocatesPhysDest = 1'b0;
    end
  end

  always @(*) begin
    if(uopNeedsNewPhysDest) begin
      io_renamedUopsOut_0_rename_physDest_idx = io_physRegsIn_0;
    end else begin
      io_renamedUopsOut_0_rename_physDest_idx = 6'h0;
    end
  end

  always @(*) begin
    if(uopNeedsNewPhysDest) begin
      io_renamedUopsOut_0_rename_physDestIsFpr = (io_decodedUopsIn_0_archDest_rtype == ArchRegType_FPR);
    end else begin
      io_renamedUopsOut_0_rename_physDestIsFpr = 1'b0;
    end
  end

  assign io_ratWritePorts_0_wen = uopNeedsNewPhysDest;
  assign io_ratWritePorts_0_archReg = io_decodedUopsIn_0_archDest_idx;
  assign io_ratWritePorts_0_physReg = io_physRegsIn_0;
  assign _zz_1 = (io_decodedUopsIn_0_archDest_rtype == ArchRegType_FPR);
  assign _zz_2 = (io_decodedUopsIn_0_archSrc1_rtype == ArchRegType_FPR);
  assign _zz_3 = (io_decodedUopsIn_0_archSrc2_rtype == ArchRegType_FPR);
  assign _zz_4 = (io_decodedUopsIn_0_archDest_rtype == ArchRegType_FPR);
  always @(posedge clk) begin
    if(reset) begin
    end else begin
      if(uopNeedsNewPhysDest) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // RenameUnit.scala:L100
          `else
            if(!1'b0) begin
              $display("NOTE(RenameUnit.scala:100):  [RenameUnit] Rename for uop@%x: archDest=%x -> physReg=%x (isFPR=%x)Src1: archSrc1=%x -> physReg=%x (isFPR=%x, bypassed=0)Src2: archSrc2=%x -> physReg=%x (isFPR=%x, bypassed=0)oldPhysDest: archDest=%x -> oldPhysReg=%x (isFPR=%x)", io_decodedUopsIn_0_pc, io_decodedUopsIn_0_archDest_idx, io_physRegsIn_0, _zz_1, io_decodedUopsIn_0_archSrc1_idx, io_renamedUopsOut_0_rename_physSrc1_idx, _zz_2, io_decodedUopsIn_0_archSrc2_idx, io_renamedUopsOut_0_rename_physSrc2_idx, _zz_3, io_decodedUopsIn_0_archDest_idx, io_renamedUopsOut_0_rename_oldPhysDest_idx, _zz_4); // RenameUnit.scala:L100
            end
          `endif
        `endif
      end
    end
  end

  always @(posedge clk) begin
    toplevel_RenamePlugin_setup_renameUnit_debugDecodedArchSrc2 <= io_decodedUopsIn_0_archSrc2_idx;
    toplevel_RenamePlugin_setup_renameUnit_debugDecodedUseArchSrc2 <= io_decodedUopsIn_0_useArchSrc2;
    toplevel_RenamePlugin_setup_renameUnit_debugRenamedPhysSrc2 <= io_renamedUopsOut_0_rename_physSrc2_idx;
  end


endmodule

//OneShot_4 replaced by OneShot

//OneShot_3 replaced by OneShot

//OneShot_2 replaced by OneShot

//OneShot_1 replaced by OneShot

module SimpleFreeList (
  input  wire          io_allocate_0_enable,
  output wire [5:0]    io_allocate_0_physReg,
  output wire          io_allocate_0_success,
  input  wire          io_free_0_enable,
  input  wire [5:0]    io_free_0_physReg,
  input  wire          io_recover,
  output wire [5:0]    io_numFreeRegs,
  input  wire          clk,
  input  wire          reset
);

  reg        [0:0]    _zz_freeCount;
  wire       [0:0]    _zz_freeCount_1;
  wire       [5:0]    _zz_availableToAlloc;
  reg        [0:0]    _zz_allocCount;
  wire       [0:0]    _zz_allocCount_1;
  wire       [4:0]    _zz__zz_1;
  wire       [4:0]    _zz__zz_io_allocate_0_physReg;
  wire       [4:0]    _zz__zz_io_allocate_0_physReg_1;
  reg        [5:0]    _zz__zz_io_allocate_0_physReg_2;
  wire       [4:0]    _zz__zz_io_allocate_0_physReg_3;
  wire       [4:0]    _zz_allocPtr;
  wire       [4:0]    _zz_freePtr;
  wire       [5:0]    _zz_occupancyCounter;
  wire       [5:0]    _zz_occupancyCounter_1;
  wire       [5:0]    _zz_occupancyCounter_2;
  reg        [5:0]    dataVec_0;
  reg        [5:0]    dataVec_1;
  reg        [5:0]    dataVec_2;
  reg        [5:0]    dataVec_3;
  reg        [5:0]    dataVec_4;
  reg        [5:0]    dataVec_5;
  reg        [5:0]    dataVec_6;
  reg        [5:0]    dataVec_7;
  reg        [5:0]    dataVec_8;
  reg        [5:0]    dataVec_9;
  reg        [5:0]    dataVec_10;
  reg        [5:0]    dataVec_11;
  reg        [5:0]    dataVec_12;
  reg        [5:0]    dataVec_13;
  reg        [5:0]    dataVec_14;
  reg        [5:0]    dataVec_15;
  reg        [5:0]    dataVec_16;
  reg        [5:0]    dataVec_17;
  reg        [5:0]    dataVec_18;
  reg        [5:0]    dataVec_19;
  reg        [5:0]    dataVec_20;
  reg        [5:0]    dataVec_21;
  reg        [5:0]    dataVec_22;
  reg        [5:0]    dataVec_23;
  reg        [5:0]    dataVec_24;
  reg        [5:0]    dataVec_25;
  reg        [5:0]    dataVec_26;
  reg        [5:0]    dataVec_27;
  reg        [5:0]    dataVec_28;
  reg        [5:0]    dataVec_29;
  reg        [5:0]    dataVec_30;
  reg        [5:0]    dataVec_31;
  reg        [4:0]    allocPtr;
  reg        [4:0]    freePtr;
  wire                isFull;
  reg        [5:0]    occupancyCounter;
  wire       [5:0]    availableToFree;
  wire                freeGrants_0;
  wire       [0:0]    freeCount;
  wire       [5:0]    availableToAlloc;
  wire                allocateGrants_0;
  wire       [0:0]    allocCount;
  wire       [31:0]   _zz_1;
  reg                 allocateGrants_0_regNext;
  reg        [5:0]    _zz_io_allocate_0_physReg;
  reg                 freeGrantsReg_0;

  assign _zz_availableToAlloc = {5'd0, freeCount};
  assign _zz__zz_1 = (freePtr + 5'h0);
  assign _zz__zz_io_allocate_0_physReg = (freePtr + 5'h0);
  assign _zz__zz_io_allocate_0_physReg_1 = (allocPtr + 5'h0);
  assign _zz__zz_io_allocate_0_physReg_3 = (allocPtr + 5'h0);
  assign _zz_allocPtr = {4'd0, allocCount};
  assign _zz_freePtr = {4'd0, freeCount};
  assign _zz_occupancyCounter = (occupancyCounter + _zz_occupancyCounter_1);
  assign _zz_occupancyCounter_1 = {5'd0, freeCount};
  assign _zz_occupancyCounter_2 = {5'd0, allocCount};
  assign _zz_freeCount_1 = freeGrants_0;
  assign _zz_allocCount_1 = allocateGrants_0;
  always @(*) begin
    case(_zz_freeCount_1)
      1'b0 : _zz_freeCount = 1'b0;
      default : _zz_freeCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_allocCount_1)
      1'b0 : _zz_allocCount = 1'b0;
      default : _zz_allocCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_allocate_0_physReg_3)
      5'b00000 : _zz__zz_io_allocate_0_physReg_2 = dataVec_0;
      5'b00001 : _zz__zz_io_allocate_0_physReg_2 = dataVec_1;
      5'b00010 : _zz__zz_io_allocate_0_physReg_2 = dataVec_2;
      5'b00011 : _zz__zz_io_allocate_0_physReg_2 = dataVec_3;
      5'b00100 : _zz__zz_io_allocate_0_physReg_2 = dataVec_4;
      5'b00101 : _zz__zz_io_allocate_0_physReg_2 = dataVec_5;
      5'b00110 : _zz__zz_io_allocate_0_physReg_2 = dataVec_6;
      5'b00111 : _zz__zz_io_allocate_0_physReg_2 = dataVec_7;
      5'b01000 : _zz__zz_io_allocate_0_physReg_2 = dataVec_8;
      5'b01001 : _zz__zz_io_allocate_0_physReg_2 = dataVec_9;
      5'b01010 : _zz__zz_io_allocate_0_physReg_2 = dataVec_10;
      5'b01011 : _zz__zz_io_allocate_0_physReg_2 = dataVec_11;
      5'b01100 : _zz__zz_io_allocate_0_physReg_2 = dataVec_12;
      5'b01101 : _zz__zz_io_allocate_0_physReg_2 = dataVec_13;
      5'b01110 : _zz__zz_io_allocate_0_physReg_2 = dataVec_14;
      5'b01111 : _zz__zz_io_allocate_0_physReg_2 = dataVec_15;
      5'b10000 : _zz__zz_io_allocate_0_physReg_2 = dataVec_16;
      5'b10001 : _zz__zz_io_allocate_0_physReg_2 = dataVec_17;
      5'b10010 : _zz__zz_io_allocate_0_physReg_2 = dataVec_18;
      5'b10011 : _zz__zz_io_allocate_0_physReg_2 = dataVec_19;
      5'b10100 : _zz__zz_io_allocate_0_physReg_2 = dataVec_20;
      5'b10101 : _zz__zz_io_allocate_0_physReg_2 = dataVec_21;
      5'b10110 : _zz__zz_io_allocate_0_physReg_2 = dataVec_22;
      5'b10111 : _zz__zz_io_allocate_0_physReg_2 = dataVec_23;
      5'b11000 : _zz__zz_io_allocate_0_physReg_2 = dataVec_24;
      5'b11001 : _zz__zz_io_allocate_0_physReg_2 = dataVec_25;
      5'b11010 : _zz__zz_io_allocate_0_physReg_2 = dataVec_26;
      5'b11011 : _zz__zz_io_allocate_0_physReg_2 = dataVec_27;
      5'b11100 : _zz__zz_io_allocate_0_physReg_2 = dataVec_28;
      5'b11101 : _zz__zz_io_allocate_0_physReg_2 = dataVec_29;
      5'b11110 : _zz__zz_io_allocate_0_physReg_2 = dataVec_30;
      default : _zz__zz_io_allocate_0_physReg_2 = dataVec_31;
    endcase
  end

  assign isFull = 1'b1;
  assign availableToFree = (6'h20 - occupancyCounter);
  assign freeGrants_0 = (((! io_recover) && io_free_0_enable) && (6'h0 < availableToFree));
  assign freeCount = _zz_freeCount;
  assign availableToAlloc = (occupancyCounter + _zz_availableToAlloc);
  assign allocateGrants_0 = (((! io_recover) && io_allocate_0_enable) && (6'h0 < availableToAlloc));
  assign allocCount = _zz_allocCount;
  assign _zz_1 = ({31'd0,1'b1} <<< _zz__zz_1);
  assign io_allocate_0_success = allocateGrants_0_regNext;
  assign io_allocate_0_physReg = _zz_io_allocate_0_physReg;
  assign io_numFreeRegs = occupancyCounter;
  always @(posedge clk) begin
    if(reset) begin
      dataVec_0 <= 6'h20;
      dataVec_1 <= 6'h21;
      dataVec_2 <= 6'h22;
      dataVec_3 <= 6'h23;
      dataVec_4 <= 6'h24;
      dataVec_5 <= 6'h25;
      dataVec_6 <= 6'h26;
      dataVec_7 <= 6'h27;
      dataVec_8 <= 6'h28;
      dataVec_9 <= 6'h29;
      dataVec_10 <= 6'h2a;
      dataVec_11 <= 6'h2b;
      dataVec_12 <= 6'h2c;
      dataVec_13 <= 6'h2d;
      dataVec_14 <= 6'h2e;
      dataVec_15 <= 6'h2f;
      dataVec_16 <= 6'h30;
      dataVec_17 <= 6'h31;
      dataVec_18 <= 6'h32;
      dataVec_19 <= 6'h33;
      dataVec_20 <= 6'h34;
      dataVec_21 <= 6'h35;
      dataVec_22 <= 6'h36;
      dataVec_23 <= 6'h37;
      dataVec_24 <= 6'h38;
      dataVec_25 <= 6'h39;
      dataVec_26 <= 6'h3a;
      dataVec_27 <= 6'h3b;
      dataVec_28 <= 6'h3c;
      dataVec_29 <= 6'h3d;
      dataVec_30 <= 6'h3e;
      dataVec_31 <= 6'h3f;
      allocPtr <= 5'h0;
      freePtr <= 5'h0;
      occupancyCounter <= 6'h20;
      allocateGrants_0_regNext <= 1'b0;
      freeGrantsReg_0 <= 1'b0;
    end else begin
      if(freeGrants_0) begin
        if(_zz_1[0]) begin
          dataVec_0 <= io_free_0_physReg;
        end
        if(_zz_1[1]) begin
          dataVec_1 <= io_free_0_physReg;
        end
        if(_zz_1[2]) begin
          dataVec_2 <= io_free_0_physReg;
        end
        if(_zz_1[3]) begin
          dataVec_3 <= io_free_0_physReg;
        end
        if(_zz_1[4]) begin
          dataVec_4 <= io_free_0_physReg;
        end
        if(_zz_1[5]) begin
          dataVec_5 <= io_free_0_physReg;
        end
        if(_zz_1[6]) begin
          dataVec_6 <= io_free_0_physReg;
        end
        if(_zz_1[7]) begin
          dataVec_7 <= io_free_0_physReg;
        end
        if(_zz_1[8]) begin
          dataVec_8 <= io_free_0_physReg;
        end
        if(_zz_1[9]) begin
          dataVec_9 <= io_free_0_physReg;
        end
        if(_zz_1[10]) begin
          dataVec_10 <= io_free_0_physReg;
        end
        if(_zz_1[11]) begin
          dataVec_11 <= io_free_0_physReg;
        end
        if(_zz_1[12]) begin
          dataVec_12 <= io_free_0_physReg;
        end
        if(_zz_1[13]) begin
          dataVec_13 <= io_free_0_physReg;
        end
        if(_zz_1[14]) begin
          dataVec_14 <= io_free_0_physReg;
        end
        if(_zz_1[15]) begin
          dataVec_15 <= io_free_0_physReg;
        end
        if(_zz_1[16]) begin
          dataVec_16 <= io_free_0_physReg;
        end
        if(_zz_1[17]) begin
          dataVec_17 <= io_free_0_physReg;
        end
        if(_zz_1[18]) begin
          dataVec_18 <= io_free_0_physReg;
        end
        if(_zz_1[19]) begin
          dataVec_19 <= io_free_0_physReg;
        end
        if(_zz_1[20]) begin
          dataVec_20 <= io_free_0_physReg;
        end
        if(_zz_1[21]) begin
          dataVec_21 <= io_free_0_physReg;
        end
        if(_zz_1[22]) begin
          dataVec_22 <= io_free_0_physReg;
        end
        if(_zz_1[23]) begin
          dataVec_23 <= io_free_0_physReg;
        end
        if(_zz_1[24]) begin
          dataVec_24 <= io_free_0_physReg;
        end
        if(_zz_1[25]) begin
          dataVec_25 <= io_free_0_physReg;
        end
        if(_zz_1[26]) begin
          dataVec_26 <= io_free_0_physReg;
        end
        if(_zz_1[27]) begin
          dataVec_27 <= io_free_0_physReg;
        end
        if(_zz_1[28]) begin
          dataVec_28 <= io_free_0_physReg;
        end
        if(_zz_1[29]) begin
          dataVec_29 <= io_free_0_physReg;
        end
        if(_zz_1[30]) begin
          dataVec_30 <= io_free_0_physReg;
        end
        if(_zz_1[31]) begin
          dataVec_31 <= io_free_0_physReg;
        end
      end
      allocateGrants_0_regNext <= allocateGrants_0;
      if(io_recover) begin
        allocPtr <= 5'h0;
        freePtr <= 5'h0;
        occupancyCounter <= 6'h20;
      end else begin
        allocPtr <= (allocPtr + _zz_allocPtr);
        freePtr <= (freePtr + _zz_freePtr);
        occupancyCounter <= (_zz_occupancyCounter - _zz_occupancyCounter_2);
      end
      freeGrantsReg_0 <= freeGrants_0;
    end
  end

  always @(posedge clk) begin
    if(allocateGrants_0) begin
      _zz_io_allocate_0_physReg <= ((freeGrants_0 && (_zz__zz_io_allocate_0_physReg == _zz__zz_io_allocate_0_physReg_1)) ? io_free_0_physReg : _zz__zz_io_allocate_0_physReg_2);
    end else begin
      _zz_io_allocate_0_physReg <= 6'h0;
    end
  end


endmodule

module RenameMapTable (
  input  wire [4:0]    io_readPorts_0_archReg,
  output reg  [5:0]    io_readPorts_0_physReg,
  input  wire [4:0]    io_readPorts_1_archReg,
  output reg  [5:0]    io_readPorts_1_physReg,
  input  wire [4:0]    io_readPorts_2_archReg,
  output reg  [5:0]    io_readPorts_2_physReg,
  input  wire          io_writePorts_0_wen,
  input  wire [4:0]    io_writePorts_0_archReg,
  input  wire [5:0]    io_writePorts_0_physReg,
  output wire [5:0]    io_currentState_mapping_0,
  output wire [5:0]    io_currentState_mapping_1,
  output wire [5:0]    io_currentState_mapping_2,
  output wire [5:0]    io_currentState_mapping_3,
  output wire [5:0]    io_currentState_mapping_4,
  output wire [5:0]    io_currentState_mapping_5,
  output wire [5:0]    io_currentState_mapping_6,
  output wire [5:0]    io_currentState_mapping_7,
  output wire [5:0]    io_currentState_mapping_8,
  output wire [5:0]    io_currentState_mapping_9,
  output wire [5:0]    io_currentState_mapping_10,
  output wire [5:0]    io_currentState_mapping_11,
  output wire [5:0]    io_currentState_mapping_12,
  output wire [5:0]    io_currentState_mapping_13,
  output wire [5:0]    io_currentState_mapping_14,
  output wire [5:0]    io_currentState_mapping_15,
  output wire [5:0]    io_currentState_mapping_16,
  output wire [5:0]    io_currentState_mapping_17,
  output wire [5:0]    io_currentState_mapping_18,
  output wire [5:0]    io_currentState_mapping_19,
  output wire [5:0]    io_currentState_mapping_20,
  output wire [5:0]    io_currentState_mapping_21,
  output wire [5:0]    io_currentState_mapping_22,
  output wire [5:0]    io_currentState_mapping_23,
  output wire [5:0]    io_currentState_mapping_24,
  output wire [5:0]    io_currentState_mapping_25,
  output wire [5:0]    io_currentState_mapping_26,
  output wire [5:0]    io_currentState_mapping_27,
  output wire [5:0]    io_currentState_mapping_28,
  output wire [5:0]    io_currentState_mapping_29,
  output wire [5:0]    io_currentState_mapping_30,
  output wire [5:0]    io_currentState_mapping_31,
  input  wire          io_checkpointRestore_valid,
  output wire          io_checkpointRestore_ready,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_0,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_1,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_2,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_3,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_4,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_5,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_6,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_7,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_8,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_9,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_10,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_11,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_12,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_13,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_14,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_15,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_16,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_17,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_18,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_19,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_20,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_21,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_22,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_23,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_24,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_25,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_26,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_27,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_28,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_29,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_30,
  input  wire [5:0]    io_checkpointRestore_payload_mapping_31,
  input  wire          io_checkpointSave_valid,
  output wire          io_checkpointSave_ready,
  input  wire [5:0]    io_checkpointSave_payload_mapping_0,
  input  wire [5:0]    io_checkpointSave_payload_mapping_1,
  input  wire [5:0]    io_checkpointSave_payload_mapping_2,
  input  wire [5:0]    io_checkpointSave_payload_mapping_3,
  input  wire [5:0]    io_checkpointSave_payload_mapping_4,
  input  wire [5:0]    io_checkpointSave_payload_mapping_5,
  input  wire [5:0]    io_checkpointSave_payload_mapping_6,
  input  wire [5:0]    io_checkpointSave_payload_mapping_7,
  input  wire [5:0]    io_checkpointSave_payload_mapping_8,
  input  wire [5:0]    io_checkpointSave_payload_mapping_9,
  input  wire [5:0]    io_checkpointSave_payload_mapping_10,
  input  wire [5:0]    io_checkpointSave_payload_mapping_11,
  input  wire [5:0]    io_checkpointSave_payload_mapping_12,
  input  wire [5:0]    io_checkpointSave_payload_mapping_13,
  input  wire [5:0]    io_checkpointSave_payload_mapping_14,
  input  wire [5:0]    io_checkpointSave_payload_mapping_15,
  input  wire [5:0]    io_checkpointSave_payload_mapping_16,
  input  wire [5:0]    io_checkpointSave_payload_mapping_17,
  input  wire [5:0]    io_checkpointSave_payload_mapping_18,
  input  wire [5:0]    io_checkpointSave_payload_mapping_19,
  input  wire [5:0]    io_checkpointSave_payload_mapping_20,
  input  wire [5:0]    io_checkpointSave_payload_mapping_21,
  input  wire [5:0]    io_checkpointSave_payload_mapping_22,
  input  wire [5:0]    io_checkpointSave_payload_mapping_23,
  input  wire [5:0]    io_checkpointSave_payload_mapping_24,
  input  wire [5:0]    io_checkpointSave_payload_mapping_25,
  input  wire [5:0]    io_checkpointSave_payload_mapping_26,
  input  wire [5:0]    io_checkpointSave_payload_mapping_27,
  input  wire [5:0]    io_checkpointSave_payload_mapping_28,
  input  wire [5:0]    io_checkpointSave_payload_mapping_29,
  input  wire [5:0]    io_checkpointSave_payload_mapping_30,
  input  wire [5:0]    io_checkpointSave_payload_mapping_31,
  input  wire          clk,
  input  wire          reset
);

  reg        [5:0]    _zz_io_readPorts_0_physReg;
  reg        [5:0]    _zz_io_readPorts_1_physReg;
  reg        [5:0]    _zz_io_readPorts_2_physReg;
  reg        [5:0]    mapReg_mapping_0;
  reg        [5:0]    mapReg_mapping_1;
  reg        [5:0]    mapReg_mapping_2;
  reg        [5:0]    mapReg_mapping_3;
  reg        [5:0]    mapReg_mapping_4;
  reg        [5:0]    mapReg_mapping_5;
  reg        [5:0]    mapReg_mapping_6;
  reg        [5:0]    mapReg_mapping_7;
  reg        [5:0]    mapReg_mapping_8;
  reg        [5:0]    mapReg_mapping_9;
  reg        [5:0]    mapReg_mapping_10;
  reg        [5:0]    mapReg_mapping_11;
  reg        [5:0]    mapReg_mapping_12;
  reg        [5:0]    mapReg_mapping_13;
  reg        [5:0]    mapReg_mapping_14;
  reg        [5:0]    mapReg_mapping_15;
  reg        [5:0]    mapReg_mapping_16;
  reg        [5:0]    mapReg_mapping_17;
  reg        [5:0]    mapReg_mapping_18;
  reg        [5:0]    mapReg_mapping_19;
  reg        [5:0]    mapReg_mapping_20;
  reg        [5:0]    mapReg_mapping_21;
  reg        [5:0]    mapReg_mapping_22;
  reg        [5:0]    mapReg_mapping_23;
  reg        [5:0]    mapReg_mapping_24;
  reg        [5:0]    mapReg_mapping_25;
  reg        [5:0]    mapReg_mapping_26;
  reg        [5:0]    mapReg_mapping_27;
  reg        [5:0]    mapReg_mapping_28;
  reg        [5:0]    mapReg_mapping_29;
  reg        [5:0]    mapReg_mapping_30;
  reg        [5:0]    mapReg_mapping_31;
  reg        [5:0]    nextMapRegMapping_0;
  reg        [5:0]    nextMapRegMapping_1;
  reg        [5:0]    nextMapRegMapping_2;
  reg        [5:0]    nextMapRegMapping_3;
  reg        [5:0]    nextMapRegMapping_4;
  reg        [5:0]    nextMapRegMapping_5;
  reg        [5:0]    nextMapRegMapping_6;
  reg        [5:0]    nextMapRegMapping_7;
  reg        [5:0]    nextMapRegMapping_8;
  reg        [5:0]    nextMapRegMapping_9;
  reg        [5:0]    nextMapRegMapping_10;
  reg        [5:0]    nextMapRegMapping_11;
  reg        [5:0]    nextMapRegMapping_12;
  reg        [5:0]    nextMapRegMapping_13;
  reg        [5:0]    nextMapRegMapping_14;
  reg        [5:0]    nextMapRegMapping_15;
  reg        [5:0]    nextMapRegMapping_16;
  reg        [5:0]    nextMapRegMapping_17;
  reg        [5:0]    nextMapRegMapping_18;
  reg        [5:0]    nextMapRegMapping_19;
  reg        [5:0]    nextMapRegMapping_20;
  reg        [5:0]    nextMapRegMapping_21;
  reg        [5:0]    nextMapRegMapping_22;
  reg        [5:0]    nextMapRegMapping_23;
  reg        [5:0]    nextMapRegMapping_24;
  reg        [5:0]    nextMapRegMapping_25;
  reg        [5:0]    nextMapRegMapping_26;
  reg        [5:0]    nextMapRegMapping_27;
  reg        [5:0]    nextMapRegMapping_28;
  reg        [5:0]    nextMapRegMapping_29;
  reg        [5:0]    nextMapRegMapping_30;
  reg        [5:0]    nextMapRegMapping_31;
  wire                when_RenameMapTable_l120;
  wire                when_RenameMapTable_l120_1;
  wire                when_RenameMapTable_l120_2;
  wire                when_RenameMapTable_l138;
  wire       [31:0]   _zz_1;

  always @(*) begin
    case(io_readPorts_0_archReg)
      5'b00000 : _zz_io_readPorts_0_physReg = mapReg_mapping_0;
      5'b00001 : _zz_io_readPorts_0_physReg = mapReg_mapping_1;
      5'b00010 : _zz_io_readPorts_0_physReg = mapReg_mapping_2;
      5'b00011 : _zz_io_readPorts_0_physReg = mapReg_mapping_3;
      5'b00100 : _zz_io_readPorts_0_physReg = mapReg_mapping_4;
      5'b00101 : _zz_io_readPorts_0_physReg = mapReg_mapping_5;
      5'b00110 : _zz_io_readPorts_0_physReg = mapReg_mapping_6;
      5'b00111 : _zz_io_readPorts_0_physReg = mapReg_mapping_7;
      5'b01000 : _zz_io_readPorts_0_physReg = mapReg_mapping_8;
      5'b01001 : _zz_io_readPorts_0_physReg = mapReg_mapping_9;
      5'b01010 : _zz_io_readPorts_0_physReg = mapReg_mapping_10;
      5'b01011 : _zz_io_readPorts_0_physReg = mapReg_mapping_11;
      5'b01100 : _zz_io_readPorts_0_physReg = mapReg_mapping_12;
      5'b01101 : _zz_io_readPorts_0_physReg = mapReg_mapping_13;
      5'b01110 : _zz_io_readPorts_0_physReg = mapReg_mapping_14;
      5'b01111 : _zz_io_readPorts_0_physReg = mapReg_mapping_15;
      5'b10000 : _zz_io_readPorts_0_physReg = mapReg_mapping_16;
      5'b10001 : _zz_io_readPorts_0_physReg = mapReg_mapping_17;
      5'b10010 : _zz_io_readPorts_0_physReg = mapReg_mapping_18;
      5'b10011 : _zz_io_readPorts_0_physReg = mapReg_mapping_19;
      5'b10100 : _zz_io_readPorts_0_physReg = mapReg_mapping_20;
      5'b10101 : _zz_io_readPorts_0_physReg = mapReg_mapping_21;
      5'b10110 : _zz_io_readPorts_0_physReg = mapReg_mapping_22;
      5'b10111 : _zz_io_readPorts_0_physReg = mapReg_mapping_23;
      5'b11000 : _zz_io_readPorts_0_physReg = mapReg_mapping_24;
      5'b11001 : _zz_io_readPorts_0_physReg = mapReg_mapping_25;
      5'b11010 : _zz_io_readPorts_0_physReg = mapReg_mapping_26;
      5'b11011 : _zz_io_readPorts_0_physReg = mapReg_mapping_27;
      5'b11100 : _zz_io_readPorts_0_physReg = mapReg_mapping_28;
      5'b11101 : _zz_io_readPorts_0_physReg = mapReg_mapping_29;
      5'b11110 : _zz_io_readPorts_0_physReg = mapReg_mapping_30;
      default : _zz_io_readPorts_0_physReg = mapReg_mapping_31;
    endcase
  end

  always @(*) begin
    case(io_readPorts_1_archReg)
      5'b00000 : _zz_io_readPorts_1_physReg = mapReg_mapping_0;
      5'b00001 : _zz_io_readPorts_1_physReg = mapReg_mapping_1;
      5'b00010 : _zz_io_readPorts_1_physReg = mapReg_mapping_2;
      5'b00011 : _zz_io_readPorts_1_physReg = mapReg_mapping_3;
      5'b00100 : _zz_io_readPorts_1_physReg = mapReg_mapping_4;
      5'b00101 : _zz_io_readPorts_1_physReg = mapReg_mapping_5;
      5'b00110 : _zz_io_readPorts_1_physReg = mapReg_mapping_6;
      5'b00111 : _zz_io_readPorts_1_physReg = mapReg_mapping_7;
      5'b01000 : _zz_io_readPorts_1_physReg = mapReg_mapping_8;
      5'b01001 : _zz_io_readPorts_1_physReg = mapReg_mapping_9;
      5'b01010 : _zz_io_readPorts_1_physReg = mapReg_mapping_10;
      5'b01011 : _zz_io_readPorts_1_physReg = mapReg_mapping_11;
      5'b01100 : _zz_io_readPorts_1_physReg = mapReg_mapping_12;
      5'b01101 : _zz_io_readPorts_1_physReg = mapReg_mapping_13;
      5'b01110 : _zz_io_readPorts_1_physReg = mapReg_mapping_14;
      5'b01111 : _zz_io_readPorts_1_physReg = mapReg_mapping_15;
      5'b10000 : _zz_io_readPorts_1_physReg = mapReg_mapping_16;
      5'b10001 : _zz_io_readPorts_1_physReg = mapReg_mapping_17;
      5'b10010 : _zz_io_readPorts_1_physReg = mapReg_mapping_18;
      5'b10011 : _zz_io_readPorts_1_physReg = mapReg_mapping_19;
      5'b10100 : _zz_io_readPorts_1_physReg = mapReg_mapping_20;
      5'b10101 : _zz_io_readPorts_1_physReg = mapReg_mapping_21;
      5'b10110 : _zz_io_readPorts_1_physReg = mapReg_mapping_22;
      5'b10111 : _zz_io_readPorts_1_physReg = mapReg_mapping_23;
      5'b11000 : _zz_io_readPorts_1_physReg = mapReg_mapping_24;
      5'b11001 : _zz_io_readPorts_1_physReg = mapReg_mapping_25;
      5'b11010 : _zz_io_readPorts_1_physReg = mapReg_mapping_26;
      5'b11011 : _zz_io_readPorts_1_physReg = mapReg_mapping_27;
      5'b11100 : _zz_io_readPorts_1_physReg = mapReg_mapping_28;
      5'b11101 : _zz_io_readPorts_1_physReg = mapReg_mapping_29;
      5'b11110 : _zz_io_readPorts_1_physReg = mapReg_mapping_30;
      default : _zz_io_readPorts_1_physReg = mapReg_mapping_31;
    endcase
  end

  always @(*) begin
    case(io_readPorts_2_archReg)
      5'b00000 : _zz_io_readPorts_2_physReg = mapReg_mapping_0;
      5'b00001 : _zz_io_readPorts_2_physReg = mapReg_mapping_1;
      5'b00010 : _zz_io_readPorts_2_physReg = mapReg_mapping_2;
      5'b00011 : _zz_io_readPorts_2_physReg = mapReg_mapping_3;
      5'b00100 : _zz_io_readPorts_2_physReg = mapReg_mapping_4;
      5'b00101 : _zz_io_readPorts_2_physReg = mapReg_mapping_5;
      5'b00110 : _zz_io_readPorts_2_physReg = mapReg_mapping_6;
      5'b00111 : _zz_io_readPorts_2_physReg = mapReg_mapping_7;
      5'b01000 : _zz_io_readPorts_2_physReg = mapReg_mapping_8;
      5'b01001 : _zz_io_readPorts_2_physReg = mapReg_mapping_9;
      5'b01010 : _zz_io_readPorts_2_physReg = mapReg_mapping_10;
      5'b01011 : _zz_io_readPorts_2_physReg = mapReg_mapping_11;
      5'b01100 : _zz_io_readPorts_2_physReg = mapReg_mapping_12;
      5'b01101 : _zz_io_readPorts_2_physReg = mapReg_mapping_13;
      5'b01110 : _zz_io_readPorts_2_physReg = mapReg_mapping_14;
      5'b01111 : _zz_io_readPorts_2_physReg = mapReg_mapping_15;
      5'b10000 : _zz_io_readPorts_2_physReg = mapReg_mapping_16;
      5'b10001 : _zz_io_readPorts_2_physReg = mapReg_mapping_17;
      5'b10010 : _zz_io_readPorts_2_physReg = mapReg_mapping_18;
      5'b10011 : _zz_io_readPorts_2_physReg = mapReg_mapping_19;
      5'b10100 : _zz_io_readPorts_2_physReg = mapReg_mapping_20;
      5'b10101 : _zz_io_readPorts_2_physReg = mapReg_mapping_21;
      5'b10110 : _zz_io_readPorts_2_physReg = mapReg_mapping_22;
      5'b10111 : _zz_io_readPorts_2_physReg = mapReg_mapping_23;
      5'b11000 : _zz_io_readPorts_2_physReg = mapReg_mapping_24;
      5'b11001 : _zz_io_readPorts_2_physReg = mapReg_mapping_25;
      5'b11010 : _zz_io_readPorts_2_physReg = mapReg_mapping_26;
      5'b11011 : _zz_io_readPorts_2_physReg = mapReg_mapping_27;
      5'b11100 : _zz_io_readPorts_2_physReg = mapReg_mapping_28;
      5'b11101 : _zz_io_readPorts_2_physReg = mapReg_mapping_29;
      5'b11110 : _zz_io_readPorts_2_physReg = mapReg_mapping_30;
      default : _zz_io_readPorts_2_physReg = mapReg_mapping_31;
    endcase
  end

  always @(*) begin
    nextMapRegMapping_0 = mapReg_mapping_0;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_0 = io_checkpointRestore_payload_mapping_0;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[0]) begin
          nextMapRegMapping_0 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_1 = mapReg_mapping_1;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_1 = io_checkpointRestore_payload_mapping_1;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[1]) begin
          nextMapRegMapping_1 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_2 = mapReg_mapping_2;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_2 = io_checkpointRestore_payload_mapping_2;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[2]) begin
          nextMapRegMapping_2 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_3 = mapReg_mapping_3;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_3 = io_checkpointRestore_payload_mapping_3;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[3]) begin
          nextMapRegMapping_3 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_4 = mapReg_mapping_4;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_4 = io_checkpointRestore_payload_mapping_4;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[4]) begin
          nextMapRegMapping_4 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_5 = mapReg_mapping_5;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_5 = io_checkpointRestore_payload_mapping_5;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[5]) begin
          nextMapRegMapping_5 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_6 = mapReg_mapping_6;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_6 = io_checkpointRestore_payload_mapping_6;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[6]) begin
          nextMapRegMapping_6 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_7 = mapReg_mapping_7;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_7 = io_checkpointRestore_payload_mapping_7;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[7]) begin
          nextMapRegMapping_7 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_8 = mapReg_mapping_8;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_8 = io_checkpointRestore_payload_mapping_8;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[8]) begin
          nextMapRegMapping_8 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_9 = mapReg_mapping_9;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_9 = io_checkpointRestore_payload_mapping_9;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[9]) begin
          nextMapRegMapping_9 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_10 = mapReg_mapping_10;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_10 = io_checkpointRestore_payload_mapping_10;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[10]) begin
          nextMapRegMapping_10 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_11 = mapReg_mapping_11;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_11 = io_checkpointRestore_payload_mapping_11;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[11]) begin
          nextMapRegMapping_11 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_12 = mapReg_mapping_12;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_12 = io_checkpointRestore_payload_mapping_12;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[12]) begin
          nextMapRegMapping_12 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_13 = mapReg_mapping_13;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_13 = io_checkpointRestore_payload_mapping_13;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[13]) begin
          nextMapRegMapping_13 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_14 = mapReg_mapping_14;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_14 = io_checkpointRestore_payload_mapping_14;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[14]) begin
          nextMapRegMapping_14 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_15 = mapReg_mapping_15;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_15 = io_checkpointRestore_payload_mapping_15;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[15]) begin
          nextMapRegMapping_15 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_16 = mapReg_mapping_16;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_16 = io_checkpointRestore_payload_mapping_16;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[16]) begin
          nextMapRegMapping_16 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_17 = mapReg_mapping_17;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_17 = io_checkpointRestore_payload_mapping_17;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[17]) begin
          nextMapRegMapping_17 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_18 = mapReg_mapping_18;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_18 = io_checkpointRestore_payload_mapping_18;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[18]) begin
          nextMapRegMapping_18 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_19 = mapReg_mapping_19;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_19 = io_checkpointRestore_payload_mapping_19;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[19]) begin
          nextMapRegMapping_19 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_20 = mapReg_mapping_20;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_20 = io_checkpointRestore_payload_mapping_20;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[20]) begin
          nextMapRegMapping_20 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_21 = mapReg_mapping_21;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_21 = io_checkpointRestore_payload_mapping_21;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[21]) begin
          nextMapRegMapping_21 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_22 = mapReg_mapping_22;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_22 = io_checkpointRestore_payload_mapping_22;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[22]) begin
          nextMapRegMapping_22 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_23 = mapReg_mapping_23;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_23 = io_checkpointRestore_payload_mapping_23;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[23]) begin
          nextMapRegMapping_23 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_24 = mapReg_mapping_24;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_24 = io_checkpointRestore_payload_mapping_24;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[24]) begin
          nextMapRegMapping_24 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_25 = mapReg_mapping_25;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_25 = io_checkpointRestore_payload_mapping_25;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[25]) begin
          nextMapRegMapping_25 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_26 = mapReg_mapping_26;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_26 = io_checkpointRestore_payload_mapping_26;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[26]) begin
          nextMapRegMapping_26 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_27 = mapReg_mapping_27;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_27 = io_checkpointRestore_payload_mapping_27;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[27]) begin
          nextMapRegMapping_27 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_28 = mapReg_mapping_28;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_28 = io_checkpointRestore_payload_mapping_28;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[28]) begin
          nextMapRegMapping_28 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_29 = mapReg_mapping_29;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_29 = io_checkpointRestore_payload_mapping_29;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[29]) begin
          nextMapRegMapping_29 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_30 = mapReg_mapping_30;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_30 = io_checkpointRestore_payload_mapping_30;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[30]) begin
          nextMapRegMapping_30 = io_writePorts_0_physReg;
        end
      end
    end
  end

  always @(*) begin
    nextMapRegMapping_31 = mapReg_mapping_31;
    if(io_checkpointRestore_valid) begin
      nextMapRegMapping_31 = io_checkpointRestore_payload_mapping_31;
    end else begin
      if(when_RenameMapTable_l138) begin
        if(_zz_1[31]) begin
          nextMapRegMapping_31 = io_writePorts_0_physReg;
        end
      end
    end
  end

  assign when_RenameMapTable_l120 = (io_readPorts_0_archReg == 5'h0);
  always @(*) begin
    if(when_RenameMapTable_l120) begin
      io_readPorts_0_physReg = 6'h0;
    end else begin
      io_readPorts_0_physReg = _zz_io_readPorts_0_physReg;
    end
  end

  assign when_RenameMapTable_l120_1 = (io_readPorts_1_archReg == 5'h0);
  always @(*) begin
    if(when_RenameMapTable_l120_1) begin
      io_readPorts_1_physReg = 6'h0;
    end else begin
      io_readPorts_1_physReg = _zz_io_readPorts_1_physReg;
    end
  end

  assign when_RenameMapTable_l120_2 = (io_readPorts_2_archReg == 5'h0);
  always @(*) begin
    if(when_RenameMapTable_l120_2) begin
      io_readPorts_2_physReg = 6'h0;
    end else begin
      io_readPorts_2_physReg = _zz_io_readPorts_2_physReg;
    end
  end

  assign when_RenameMapTable_l138 = (io_writePorts_0_wen && (io_writePorts_0_archReg != 5'h0));
  assign _zz_1 = ({31'd0,1'b1} <<< io_writePorts_0_archReg);
  assign io_checkpointRestore_ready = 1'b1;
  assign io_checkpointSave_ready = 1'b1;
  assign io_currentState_mapping_0 = mapReg_mapping_0;
  assign io_currentState_mapping_1 = mapReg_mapping_1;
  assign io_currentState_mapping_2 = mapReg_mapping_2;
  assign io_currentState_mapping_3 = mapReg_mapping_3;
  assign io_currentState_mapping_4 = mapReg_mapping_4;
  assign io_currentState_mapping_5 = mapReg_mapping_5;
  assign io_currentState_mapping_6 = mapReg_mapping_6;
  assign io_currentState_mapping_7 = mapReg_mapping_7;
  assign io_currentState_mapping_8 = mapReg_mapping_8;
  assign io_currentState_mapping_9 = mapReg_mapping_9;
  assign io_currentState_mapping_10 = mapReg_mapping_10;
  assign io_currentState_mapping_11 = mapReg_mapping_11;
  assign io_currentState_mapping_12 = mapReg_mapping_12;
  assign io_currentState_mapping_13 = mapReg_mapping_13;
  assign io_currentState_mapping_14 = mapReg_mapping_14;
  assign io_currentState_mapping_15 = mapReg_mapping_15;
  assign io_currentState_mapping_16 = mapReg_mapping_16;
  assign io_currentState_mapping_17 = mapReg_mapping_17;
  assign io_currentState_mapping_18 = mapReg_mapping_18;
  assign io_currentState_mapping_19 = mapReg_mapping_19;
  assign io_currentState_mapping_20 = mapReg_mapping_20;
  assign io_currentState_mapping_21 = mapReg_mapping_21;
  assign io_currentState_mapping_22 = mapReg_mapping_22;
  assign io_currentState_mapping_23 = mapReg_mapping_23;
  assign io_currentState_mapping_24 = mapReg_mapping_24;
  assign io_currentState_mapping_25 = mapReg_mapping_25;
  assign io_currentState_mapping_26 = mapReg_mapping_26;
  assign io_currentState_mapping_27 = mapReg_mapping_27;
  assign io_currentState_mapping_28 = mapReg_mapping_28;
  assign io_currentState_mapping_29 = mapReg_mapping_29;
  assign io_currentState_mapping_30 = mapReg_mapping_30;
  assign io_currentState_mapping_31 = mapReg_mapping_31;
  always @(posedge clk) begin
    if(reset) begin
      mapReg_mapping_0 <= 6'h0;
      mapReg_mapping_1 <= 6'h01;
      mapReg_mapping_2 <= 6'h02;
      mapReg_mapping_3 <= 6'h03;
      mapReg_mapping_4 <= 6'h04;
      mapReg_mapping_5 <= 6'h05;
      mapReg_mapping_6 <= 6'h06;
      mapReg_mapping_7 <= 6'h07;
      mapReg_mapping_8 <= 6'h08;
      mapReg_mapping_9 <= 6'h09;
      mapReg_mapping_10 <= 6'h0a;
      mapReg_mapping_11 <= 6'h0b;
      mapReg_mapping_12 <= 6'h0c;
      mapReg_mapping_13 <= 6'h0d;
      mapReg_mapping_14 <= 6'h0e;
      mapReg_mapping_15 <= 6'h0f;
      mapReg_mapping_16 <= 6'h10;
      mapReg_mapping_17 <= 6'h11;
      mapReg_mapping_18 <= 6'h12;
      mapReg_mapping_19 <= 6'h13;
      mapReg_mapping_20 <= 6'h14;
      mapReg_mapping_21 <= 6'h15;
      mapReg_mapping_22 <= 6'h16;
      mapReg_mapping_23 <= 6'h17;
      mapReg_mapping_24 <= 6'h18;
      mapReg_mapping_25 <= 6'h19;
      mapReg_mapping_26 <= 6'h1a;
      mapReg_mapping_27 <= 6'h1b;
      mapReg_mapping_28 <= 6'h1c;
      mapReg_mapping_29 <= 6'h1d;
      mapReg_mapping_30 <= 6'h1e;
      mapReg_mapping_31 <= 6'h1f;
    end else begin
      mapReg_mapping_0 <= nextMapRegMapping_0;
      mapReg_mapping_1 <= nextMapRegMapping_1;
      mapReg_mapping_2 <= nextMapRegMapping_2;
      mapReg_mapping_3 <= nextMapRegMapping_3;
      mapReg_mapping_4 <= nextMapRegMapping_4;
      mapReg_mapping_5 <= nextMapRegMapping_5;
      mapReg_mapping_6 <= nextMapRegMapping_6;
      mapReg_mapping_7 <= nextMapRegMapping_7;
      mapReg_mapping_8 <= nextMapRegMapping_8;
      mapReg_mapping_9 <= nextMapRegMapping_9;
      mapReg_mapping_10 <= nextMapRegMapping_10;
      mapReg_mapping_11 <= nextMapRegMapping_11;
      mapReg_mapping_12 <= nextMapRegMapping_12;
      mapReg_mapping_13 <= nextMapRegMapping_13;
      mapReg_mapping_14 <= nextMapRegMapping_14;
      mapReg_mapping_15 <= nextMapRegMapping_15;
      mapReg_mapping_16 <= nextMapRegMapping_16;
      mapReg_mapping_17 <= nextMapRegMapping_17;
      mapReg_mapping_18 <= nextMapRegMapping_18;
      mapReg_mapping_19 <= nextMapRegMapping_19;
      mapReg_mapping_20 <= nextMapRegMapping_20;
      mapReg_mapping_21 <= nextMapRegMapping_21;
      mapReg_mapping_22 <= nextMapRegMapping_22;
      mapReg_mapping_23 <= nextMapRegMapping_23;
      mapReg_mapping_24 <= nextMapRegMapping_24;
      mapReg_mapping_25 <= nextMapRegMapping_25;
      mapReg_mapping_26 <= nextMapRegMapping_26;
      mapReg_mapping_27 <= nextMapRegMapping_27;
      mapReg_mapping_28 <= nextMapRegMapping_28;
      mapReg_mapping_29 <= nextMapRegMapping_29;
      mapReg_mapping_30 <= nextMapRegMapping_30;
      mapReg_mapping_31 <= nextMapRegMapping_31;
    end
  end


endmodule

module ReorderBuffer (
  input  wire          io_allocate_0_valid,
  input  wire [31:0]   io_allocate_0_uopIn_decoded_pc,
  input  wire          io_allocate_0_uopIn_decoded_isValid,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_uopCode,
  input  wire [3:0]    io_allocate_0_uopIn_decoded_exeUnit,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_isa,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_archDest_idx,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_archDest_rtype,
  input  wire          io_allocate_0_uopIn_decoded_writeArchDestEn,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_archSrc1_idx,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_archSrc1_rtype,
  input  wire          io_allocate_0_uopIn_decoded_useArchSrc1,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_archSrc2_idx,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_archSrc2_rtype,
  input  wire          io_allocate_0_uopIn_decoded_useArchSrc2,
  input  wire          io_allocate_0_uopIn_decoded_usePcForAddr,
  input  wire [31:0]   io_allocate_0_uopIn_decoded_imm,
  input  wire [2:0]    io_allocate_0_uopIn_decoded_immUsage,
  input  wire          io_allocate_0_uopIn_decoded_aluCtrl_valid,
  input  wire          io_allocate_0_uopIn_decoded_aluCtrl_isSub,
  input  wire          io_allocate_0_uopIn_decoded_aluCtrl_isAdd,
  input  wire          io_allocate_0_uopIn_decoded_aluCtrl_isSigned,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_aluCtrl_logicOp,
  input  wire          io_allocate_0_uopIn_decoded_shiftCtrl_valid,
  input  wire          io_allocate_0_uopIn_decoded_shiftCtrl_isRight,
  input  wire          io_allocate_0_uopIn_decoded_shiftCtrl_isArithmetic,
  input  wire          io_allocate_0_uopIn_decoded_shiftCtrl_isRotate,
  input  wire          io_allocate_0_uopIn_decoded_shiftCtrl_isDoubleWord,
  input  wire          io_allocate_0_uopIn_decoded_mulDivCtrl_valid,
  input  wire          io_allocate_0_uopIn_decoded_mulDivCtrl_isDiv,
  input  wire          io_allocate_0_uopIn_decoded_mulDivCtrl_isSigned,
  input  wire          io_allocate_0_uopIn_decoded_mulDivCtrl_isWordOp,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_memCtrl_size,
  input  wire          io_allocate_0_uopIn_decoded_memCtrl_isSignedLoad,
  input  wire          io_allocate_0_uopIn_decoded_memCtrl_isStore,
  input  wire          io_allocate_0_uopIn_decoded_memCtrl_isLoadLinked,
  input  wire          io_allocate_0_uopIn_decoded_memCtrl_isStoreCond,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_memCtrl_atomicOp,
  input  wire          io_allocate_0_uopIn_decoded_memCtrl_isFence,
  input  wire [7:0]    io_allocate_0_uopIn_decoded_memCtrl_fenceMode,
  input  wire          io_allocate_0_uopIn_decoded_memCtrl_isCacheOp,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_memCtrl_cacheOpType,
  input  wire          io_allocate_0_uopIn_decoded_memCtrl_isPrefetch,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_branchCtrl_condition,
  input  wire          io_allocate_0_uopIn_decoded_branchCtrl_isJump,
  input  wire          io_allocate_0_uopIn_decoded_branchCtrl_isLink,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_branchCtrl_linkReg_idx,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype,
  input  wire          io_allocate_0_uopIn_decoded_branchCtrl_isIndirect,
  input  wire [2:0]    io_allocate_0_uopIn_decoded_branchCtrl_laCfIdx,
  input  wire [3:0]    io_allocate_0_uopIn_decoded_fpuCtrl_opType,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest,
  input  wire [2:0]    io_allocate_0_uopIn_decoded_fpuCtrl_roundingMode,
  input  wire          io_allocate_0_uopIn_decoded_fpuCtrl_isIntegerDest,
  input  wire          io_allocate_0_uopIn_decoded_fpuCtrl_isSignedCvt,
  input  wire          io_allocate_0_uopIn_decoded_fpuCtrl_fmaNegSrc1,
  input  wire [4:0]    io_allocate_0_uopIn_decoded_fpuCtrl_fcmpCond,
  input  wire [13:0]   io_allocate_0_uopIn_decoded_csrCtrl_csrAddr,
  input  wire          io_allocate_0_uopIn_decoded_csrCtrl_isWrite,
  input  wire          io_allocate_0_uopIn_decoded_csrCtrl_isRead,
  input  wire          io_allocate_0_uopIn_decoded_csrCtrl_isExchange,
  input  wire          io_allocate_0_uopIn_decoded_csrCtrl_useUimmAsSrc,
  input  wire [19:0]   io_allocate_0_uopIn_decoded_sysCtrl_sysCode,
  input  wire          io_allocate_0_uopIn_decoded_sysCtrl_isExceptionReturn,
  input  wire          io_allocate_0_uopIn_decoded_sysCtrl_isTlbOp,
  input  wire [3:0]    io_allocate_0_uopIn_decoded_sysCtrl_tlbOpType,
  input  wire [1:0]    io_allocate_0_uopIn_decoded_decodeExceptionCode,
  input  wire          io_allocate_0_uopIn_decoded_hasDecodeException,
  input  wire          io_allocate_0_uopIn_decoded_isMicrocode,
  input  wire [7:0]    io_allocate_0_uopIn_decoded_microcodeEntry,
  input  wire          io_allocate_0_uopIn_decoded_isSerializing,
  input  wire          io_allocate_0_uopIn_decoded_isBranchOrJump,
  input  wire          io_allocate_0_uopIn_decoded_branchPrediction_isTaken,
  input  wire [31:0]   io_allocate_0_uopIn_decoded_branchPrediction_target,
  input  wire          io_allocate_0_uopIn_decoded_branchPrediction_wasPredicted,
  input  wire [5:0]    io_allocate_0_uopIn_rename_physSrc1_idx,
  input  wire          io_allocate_0_uopIn_rename_physSrc1IsFpr,
  input  wire [5:0]    io_allocate_0_uopIn_rename_physSrc2_idx,
  input  wire          io_allocate_0_uopIn_rename_physSrc2IsFpr,
  input  wire [5:0]    io_allocate_0_uopIn_rename_physDest_idx,
  input  wire          io_allocate_0_uopIn_rename_physDestIsFpr,
  input  wire [5:0]    io_allocate_0_uopIn_rename_oldPhysDest_idx,
  input  wire          io_allocate_0_uopIn_rename_oldPhysDestIsFpr,
  input  wire          io_allocate_0_uopIn_rename_allocatesPhysDest,
  input  wire          io_allocate_0_uopIn_rename_writesToPhysReg,
  input  wire [3:0]    io_allocate_0_uopIn_robPtr,
  input  wire [15:0]   io_allocate_0_uopIn_uniqueId,
  input  wire          io_allocate_0_uopIn_dispatched,
  input  wire          io_allocate_0_uopIn_executed,
  input  wire          io_allocate_0_uopIn_hasException,
  input  wire [7:0]    io_allocate_0_uopIn_exceptionCode,
  input  wire [31:0]   io_allocate_0_pcIn,
  output wire [3:0]    io_allocate_0_robPtr,
  output wire          io_allocate_0_ready,
  output wire          io_canAllocate_0,
  input  wire          io_writeback_0_fire,
  input  wire [3:0]    io_writeback_0_robPtr,
  input  wire          io_writeback_0_isTaken,
  input  wire          io_writeback_0_isMispredictedBranch,
  input  wire [31:0]   io_writeback_0_result,
  input  wire          io_writeback_0_exceptionOccurred,
  input  wire [7:0]    io_writeback_0_exceptionCodeIn,
  input  wire          io_writeback_1_fire,
  input  wire [3:0]    io_writeback_1_robPtr,
  input  wire          io_writeback_1_isTaken,
  input  wire          io_writeback_1_isMispredictedBranch,
  input  wire [31:0]   io_writeback_1_result,
  input  wire          io_writeback_1_exceptionOccurred,
  input  wire [7:0]    io_writeback_1_exceptionCodeIn,
  input  wire          io_writeback_2_fire,
  input  wire [3:0]    io_writeback_2_robPtr,
  input  wire          io_writeback_2_isTaken,
  input  wire          io_writeback_2_isMispredictedBranch,
  input  wire [31:0]   io_writeback_2_result,
  input  wire          io_writeback_2_exceptionOccurred,
  input  wire [7:0]    io_writeback_2_exceptionCodeIn,
  input  wire          io_writeback_3_fire,
  input  wire [3:0]    io_writeback_3_robPtr,
  input  wire          io_writeback_3_isTaken,
  input  wire          io_writeback_3_isMispredictedBranch,
  input  wire [31:0]   io_writeback_3_result,
  input  wire          io_writeback_3_exceptionOccurred,
  input  wire [7:0]    io_writeback_3_exceptionCodeIn,
  input  wire          io_writeback_4_fire,
  input  wire [3:0]    io_writeback_4_robPtr,
  input  wire          io_writeback_4_isTaken,
  input  wire          io_writeback_4_isMispredictedBranch,
  input  wire [31:0]   io_writeback_4_result,
  input  wire          io_writeback_4_exceptionOccurred,
  input  wire [7:0]    io_writeback_4_exceptionCodeIn,
  output wire          io_commit_0_valid,
  output wire          io_commit_0_canCommit,
  output wire [31:0]   io_commit_0_entry_payload_uop_decoded_pc,
  output wire          io_commit_0_entry_payload_uop_decoded_isValid,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_uopCode,
  output wire [3:0]    io_commit_0_entry_payload_uop_decoded_exeUnit,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_isa,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_archDest_idx,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_archDest_rtype,
  output wire          io_commit_0_entry_payload_uop_decoded_writeArchDestEn,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_archSrc1_idx,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_archSrc1_rtype,
  output wire          io_commit_0_entry_payload_uop_decoded_useArchSrc1,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_archSrc2_idx,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_archSrc2_rtype,
  output wire          io_commit_0_entry_payload_uop_decoded_useArchSrc2,
  output wire          io_commit_0_entry_payload_uop_decoded_usePcForAddr,
  output wire [31:0]   io_commit_0_entry_payload_uop_decoded_imm,
  output wire [2:0]    io_commit_0_entry_payload_uop_decoded_immUsage,
  output wire          io_commit_0_entry_payload_uop_decoded_aluCtrl_valid,
  output wire          io_commit_0_entry_payload_uop_decoded_aluCtrl_isSub,
  output wire          io_commit_0_entry_payload_uop_decoded_aluCtrl_isAdd,
  output wire          io_commit_0_entry_payload_uop_decoded_aluCtrl_isSigned,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp,
  output wire          io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid,
  output wire          io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRight,
  output wire          io_commit_0_entry_payload_uop_decoded_shiftCtrl_isArithmetic,
  output wire          io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRotate,
  output wire          io_commit_0_entry_payload_uop_decoded_shiftCtrl_isDoubleWord,
  output wire          io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid,
  output wire          io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isDiv,
  output wire          io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isSigned,
  output wire          io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isWordOp,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_memCtrl_size,
  output wire          io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad,
  output wire          io_commit_0_entry_payload_uop_decoded_memCtrl_isStore,
  output wire          io_commit_0_entry_payload_uop_decoded_memCtrl_isLoadLinked,
  output wire          io_commit_0_entry_payload_uop_decoded_memCtrl_isStoreCond,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_memCtrl_atomicOp,
  output wire          io_commit_0_entry_payload_uop_decoded_memCtrl_isFence,
  output wire [7:0]    io_commit_0_entry_payload_uop_decoded_memCtrl_fenceMode,
  output wire          io_commit_0_entry_payload_uop_decoded_memCtrl_isCacheOp,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_memCtrl_cacheOpType,
  output wire          io_commit_0_entry_payload_uop_decoded_memCtrl_isPrefetch,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_branchCtrl_condition,
  output wire          io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump,
  output wire          io_commit_0_entry_payload_uop_decoded_branchCtrl_isLink,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype,
  output wire          io_commit_0_entry_payload_uop_decoded_branchCtrl_isIndirect,
  output wire [2:0]    io_commit_0_entry_payload_uop_decoded_branchCtrl_laCfIdx,
  output wire [3:0]    io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest,
  output wire [2:0]    io_commit_0_entry_payload_uop_decoded_fpuCtrl_roundingMode,
  output wire          io_commit_0_entry_payload_uop_decoded_fpuCtrl_isIntegerDest,
  output wire          io_commit_0_entry_payload_uop_decoded_fpuCtrl_isSignedCvt,
  output wire          io_commit_0_entry_payload_uop_decoded_fpuCtrl_fmaNegSrc1,
  output wire [4:0]    io_commit_0_entry_payload_uop_decoded_fpuCtrl_fcmpCond,
  output wire [13:0]   io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr,
  output wire          io_commit_0_entry_payload_uop_decoded_csrCtrl_isWrite,
  output wire          io_commit_0_entry_payload_uop_decoded_csrCtrl_isRead,
  output wire          io_commit_0_entry_payload_uop_decoded_csrCtrl_isExchange,
  output wire          io_commit_0_entry_payload_uop_decoded_csrCtrl_useUimmAsSrc,
  output wire [19:0]   io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode,
  output wire          io_commit_0_entry_payload_uop_decoded_sysCtrl_isExceptionReturn,
  output wire          io_commit_0_entry_payload_uop_decoded_sysCtrl_isTlbOp,
  output wire [3:0]    io_commit_0_entry_payload_uop_decoded_sysCtrl_tlbOpType,
  output wire [1:0]    io_commit_0_entry_payload_uop_decoded_decodeExceptionCode,
  output wire          io_commit_0_entry_payload_uop_decoded_hasDecodeException,
  output wire          io_commit_0_entry_payload_uop_decoded_isMicrocode,
  output wire [7:0]    io_commit_0_entry_payload_uop_decoded_microcodeEntry,
  output wire          io_commit_0_entry_payload_uop_decoded_isSerializing,
  output wire          io_commit_0_entry_payload_uop_decoded_isBranchOrJump,
  output wire          io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken,
  output wire [31:0]   io_commit_0_entry_payload_uop_decoded_branchPrediction_target,
  output wire          io_commit_0_entry_payload_uop_decoded_branchPrediction_wasPredicted,
  output wire [5:0]    io_commit_0_entry_payload_uop_rename_physSrc1_idx,
  output wire          io_commit_0_entry_payload_uop_rename_physSrc1IsFpr,
  output wire [5:0]    io_commit_0_entry_payload_uop_rename_physSrc2_idx,
  output wire          io_commit_0_entry_payload_uop_rename_physSrc2IsFpr,
  output wire [5:0]    io_commit_0_entry_payload_uop_rename_physDest_idx,
  output wire          io_commit_0_entry_payload_uop_rename_physDestIsFpr,
  output wire [5:0]    io_commit_0_entry_payload_uop_rename_oldPhysDest_idx,
  output wire          io_commit_0_entry_payload_uop_rename_oldPhysDestIsFpr,
  output wire          io_commit_0_entry_payload_uop_rename_allocatesPhysDest,
  output wire          io_commit_0_entry_payload_uop_rename_writesToPhysReg,
  output wire [3:0]    io_commit_0_entry_payload_uop_robPtr,
  output wire [15:0]   io_commit_0_entry_payload_uop_uniqueId,
  output wire          io_commit_0_entry_payload_uop_dispatched,
  output wire          io_commit_0_entry_payload_uop_executed,
  output wire          io_commit_0_entry_payload_uop_hasException,
  output wire [7:0]    io_commit_0_entry_payload_uop_exceptionCode,
  output wire [31:0]   io_commit_0_entry_payload_pc,
  output wire          io_commit_0_entry_status_busy,
  output wire          io_commit_0_entry_status_done,
  output wire          io_commit_0_entry_status_isMispredictedBranch,
  output wire          io_commit_0_entry_status_isTaken,
  output wire [31:0]   io_commit_0_entry_status_result,
  output wire          io_commit_0_entry_status_hasException,
  output wire [7:0]    io_commit_0_entry_status_exceptionCode,
  output wire          io_commit_0_entry_status_genBit,
  input  wire          io_commitAck_0,
  input  wire          io_flush_valid,
  input  wire [1:0]    io_flush_payload_reason,
  input  wire [3:0]    io_flush_payload_targetRobPtr,
  output reg           io_flushed,
  output wire          io_empty,
  output wire [3:0]    io_headPtrOut,
  output wire [3:0]    io_tailPtrOut,
  output wire [3:0]    io_countOut,
  input  wire          clk,
  input  wire          reset
);
  localparam BaseUopCode_NOP = 5'd0;
  localparam BaseUopCode_ILLEGAL = 5'd1;
  localparam BaseUopCode_ALU = 5'd2;
  localparam BaseUopCode_SHIFT = 5'd3;
  localparam BaseUopCode_MUL = 5'd4;
  localparam BaseUopCode_DIV = 5'd5;
  localparam BaseUopCode_LOAD = 5'd6;
  localparam BaseUopCode_STORE = 5'd7;
  localparam BaseUopCode_ATOMIC = 5'd8;
  localparam BaseUopCode_MEM_BARRIER = 5'd9;
  localparam BaseUopCode_PREFETCH = 5'd10;
  localparam BaseUopCode_BRANCH = 5'd11;
  localparam BaseUopCode_JUMP_REG = 5'd12;
  localparam BaseUopCode_JUMP_IMM = 5'd13;
  localparam BaseUopCode_SYSTEM_OP = 5'd14;
  localparam BaseUopCode_CSR_ACCESS = 5'd15;
  localparam BaseUopCode_FPU_ALU = 5'd16;
  localparam BaseUopCode_FPU_CVT = 5'd17;
  localparam BaseUopCode_FPU_CMP = 5'd18;
  localparam BaseUopCode_FPU_SEL = 5'd19;
  localparam BaseUopCode_LA_BITMANIP = 5'd20;
  localparam BaseUopCode_LA_CACOP = 5'd21;
  localparam BaseUopCode_LA_TLB = 5'd22;
  localparam BaseUopCode_IDLE = 5'd23;
  localparam ExeUnitType_NONE = 4'd0;
  localparam ExeUnitType_ALU_INT = 4'd1;
  localparam ExeUnitType_MUL_INT = 4'd2;
  localparam ExeUnitType_DIV_INT = 4'd3;
  localparam ExeUnitType_MEM = 4'd4;
  localparam ExeUnitType_BRU = 4'd5;
  localparam ExeUnitType_CSR = 4'd6;
  localparam ExeUnitType_FPU_ADD_MUL_CVT_CMP = 4'd7;
  localparam ExeUnitType_FPU_DIV_SQRT = 4'd8;
  localparam IsaType_UNKNOWN = 2'd0;
  localparam IsaType_DEMO = 2'd1;
  localparam IsaType_RISCV = 2'd2;
  localparam IsaType_LOONGARCH = 2'd3;
  localparam ArchRegType_GPR = 2'd0;
  localparam ArchRegType_FPR = 2'd1;
  localparam ArchRegType_CSR = 2'd2;
  localparam ArchRegType_LA_CF = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam MemAccessSize_B = 2'd0;
  localparam MemAccessSize_H = 2'd1;
  localparam MemAccessSize_W = 2'd2;
  localparam MemAccessSize_D = 2'd3;
  localparam BranchCondition_NUL = 5'd0;
  localparam BranchCondition_EQ = 5'd1;
  localparam BranchCondition_NE = 5'd2;
  localparam BranchCondition_LT = 5'd3;
  localparam BranchCondition_GE = 5'd4;
  localparam BranchCondition_LTU = 5'd5;
  localparam BranchCondition_GEU = 5'd6;
  localparam BranchCondition_EQZ = 5'd7;
  localparam BranchCondition_NEZ = 5'd8;
  localparam BranchCondition_LTZ = 5'd9;
  localparam BranchCondition_GEZ = 5'd10;
  localparam BranchCondition_GTZ = 5'd11;
  localparam BranchCondition_LEZ = 5'd12;
  localparam BranchCondition_F_EQ = 5'd13;
  localparam BranchCondition_F_NE = 5'd14;
  localparam BranchCondition_F_LT = 5'd15;
  localparam BranchCondition_F_LE = 5'd16;
  localparam BranchCondition_F_UN = 5'd17;
  localparam BranchCondition_LA_CF_TRUE = 5'd18;
  localparam BranchCondition_LA_CF_FALSE = 5'd19;
  localparam DecodeExCode_INVALID = 2'd0;
  localparam DecodeExCode_FETCH_ERROR = 2'd1;
  localparam DecodeExCode_DECODE_ERROR = 2'd2;
  localparam DecodeExCode_OK = 2'd3;
  localparam FlushReason_NONE = 2'd0;
  localparam FlushReason_FULL_FLUSH = 2'd1;
  localparam FlushReason_ROLLBACK_TO_ROB_IDX = 2'd2;

  wire       [369:0]  payloads_spinal_port0;
  wire       [3:0]    _zz__zz_io_allocate_0_ready;
  reg        [0:0]    _zz_numActuallyAllocatedThisCycle;
  wire       [0:0]    _zz_numActuallyAllocatedThisCycle_1;
  reg                 _zz__zz_io_commit_0_entry_status_done;
  reg                 _zz__zz_io_commit_0_entry_status_genBit;
  wire       [5:0]    _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx_1;
  wire       [5:0]    _zz_io_commit_0_entry_payload_uop_rename_physSrc2_idx;
  wire       [5:0]    _zz_io_commit_0_entry_payload_uop_rename_physDest_idx;
  wire       [5:0]    _zz_io_commit_0_entry_payload_uop_rename_oldPhysDest_idx;
  reg                 _zz_io_commit_0_entry_status_busy_1;
  reg                 _zz_io_commit_0_entry_status_isMispredictedBranch;
  reg                 _zz_io_commit_0_entry_status_isTaken;
  reg        [31:0]   _zz_io_commit_0_entry_status_result;
  reg                 _zz_io_commit_0_entry_status_hasException;
  reg        [7:0]    _zz_io_commit_0_entry_status_exceptionCode;
  reg        [0:0]    _zz_numToCommit;
  wire       [0:0]    _zz_numToCommit_1;
  wire       [3:0]    _zz_nextHead;
  wire       [3:0]    _zz_nextTail;
  wire       [3:0]    _zz_nextCount_1;
  wire       [3:0]    _zz_nextCount_2;
  wire       [3:0]    _zz_nextCount_3;
  wire       [4:0]    _zz__zz_nextCount;
  wire       [4:0]    _zz__zz_nextCount_1;
  wire       [369:0]  _zz_payloads_port;
  reg                 _zz_when_ReorderBuffer_l375_5;
  reg        [7:0]    _zz__zz_statuses_0_exceptionCode;
  reg                 _zz_when_ReorderBuffer_l375_1_1;
  reg        [7:0]    _zz__zz_statuses_0_exceptionCode_1;
  reg                 _zz_when_ReorderBuffer_l375_2_1;
  reg        [7:0]    _zz__zz_statuses_0_exceptionCode_2;
  reg                 _zz_when_ReorderBuffer_l375_3_1;
  reg        [7:0]    _zz__zz_statuses_0_exceptionCode_3;
  reg                 _zz_when_ReorderBuffer_l375_4_1;
  reg        [7:0]    _zz__zz_statuses_0_exceptionCode_4;
  wire       [3:0]    _zz__zz_when_ReorderBuffer_l418_3;
  reg                 _zz__zz_when_ReorderBuffer_l418_3_1;
  wire       [3:0]    _zz__zz_when_ReorderBuffer_l418_7;
  reg                 _zz__zz_when_ReorderBuffer_l418_7_1;
  wire       [3:0]    _zz__zz_when_ReorderBuffer_l418_11;
  reg                 _zz__zz_when_ReorderBuffer_l418_11_1;
  wire       [3:0]    _zz__zz_when_ReorderBuffer_l418_15;
  reg                 _zz__zz_when_ReorderBuffer_l418_15_1;
  wire       [3:0]    _zz__zz_when_ReorderBuffer_l418_19;
  reg                 _zz__zz_when_ReorderBuffer_l418_19_1;
  wire       [3:0]    _zz__zz_when_ReorderBuffer_l418_23;
  reg                 _zz__zz_when_ReorderBuffer_l418_23_1;
  wire       [3:0]    _zz__zz_when_ReorderBuffer_l418_27;
  reg                 _zz__zz_when_ReorderBuffer_l418_27_1;
  wire       [3:0]    _zz__zz_when_ReorderBuffer_l418_31;
  reg                 _zz__zz_when_ReorderBuffer_l418_31_1;
  reg                 _zz_1;
  reg                 statuses_0_busy;
  reg                 statuses_0_done;
  reg                 statuses_0_isMispredictedBranch;
  reg                 statuses_0_isTaken;
  reg        [31:0]   statuses_0_result;
  reg                 statuses_0_hasException;
  reg        [7:0]    statuses_0_exceptionCode;
  reg                 statuses_0_genBit;
  reg                 statuses_1_busy;
  reg                 statuses_1_done;
  reg                 statuses_1_isMispredictedBranch;
  reg                 statuses_1_isTaken;
  reg        [31:0]   statuses_1_result;
  reg                 statuses_1_hasException;
  reg        [7:0]    statuses_1_exceptionCode;
  reg                 statuses_1_genBit;
  reg                 statuses_2_busy;
  reg                 statuses_2_done;
  reg                 statuses_2_isMispredictedBranch;
  reg                 statuses_2_isTaken;
  reg        [31:0]   statuses_2_result;
  reg                 statuses_2_hasException;
  reg        [7:0]    statuses_2_exceptionCode;
  reg                 statuses_2_genBit;
  reg                 statuses_3_busy;
  reg                 statuses_3_done;
  reg                 statuses_3_isMispredictedBranch;
  reg                 statuses_3_isTaken;
  reg        [31:0]   statuses_3_result;
  reg                 statuses_3_hasException;
  reg        [7:0]    statuses_3_exceptionCode;
  reg                 statuses_3_genBit;
  reg                 statuses_4_busy;
  reg                 statuses_4_done;
  reg                 statuses_4_isMispredictedBranch;
  reg                 statuses_4_isTaken;
  reg        [31:0]   statuses_4_result;
  reg                 statuses_4_hasException;
  reg        [7:0]    statuses_4_exceptionCode;
  reg                 statuses_4_genBit;
  reg                 statuses_5_busy;
  reg                 statuses_5_done;
  reg                 statuses_5_isMispredictedBranch;
  reg                 statuses_5_isTaken;
  reg        [31:0]   statuses_5_result;
  reg                 statuses_5_hasException;
  reg        [7:0]    statuses_5_exceptionCode;
  reg                 statuses_5_genBit;
  reg                 statuses_6_busy;
  reg                 statuses_6_done;
  reg                 statuses_6_isMispredictedBranch;
  reg                 statuses_6_isTaken;
  reg        [31:0]   statuses_6_result;
  reg                 statuses_6_hasException;
  reg        [7:0]    statuses_6_exceptionCode;
  reg                 statuses_6_genBit;
  reg                 statuses_7_busy;
  reg                 statuses_7_done;
  reg                 statuses_7_isMispredictedBranch;
  reg                 statuses_7_isTaken;
  reg        [31:0]   statuses_7_result;
  reg                 statuses_7_hasException;
  reg        [7:0]    statuses_7_exceptionCode;
  reg                 statuses_7_genBit;
  reg        [3:0]    headPtr_reg;
  reg        [3:0]    tailPtr_reg;
  reg        [3:0]    count_reg;
  wire                slotWillAllocate_0;
  wire                _zz_io_allocate_0_ready;
  wire       [0:0]    numActuallyAllocatedThisCycle;
  reg                 flushInProgressReg;
  reg                 flushWasActiveLastCycle;
  wire                canCommitFlags_0;
  wire                actualCommittedMask_0;
  wire       [3:0]    _zz_canCommitFlags_0;
  wire       [2:0]    _zz_io_commit_0_entry_status_busy;
  wire                _zz_io_commit_0_entry_status_done;
  wire                _zz_io_commit_0_entry_status_genBit;
  wire       [4:0]    _zz_io_commit_0_entry_payload_uop_decoded_uopCode;
  wire       [3:0]    _zz_io_commit_0_entry_payload_uop_decoded_exeUnit;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_isa;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype;
  wire       [2:0]    _zz_io_commit_0_entry_payload_uop_decoded_immUsage;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size;
  wire       [4:0]    _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode;
  wire       [369:0]  _zz_io_commit_0_entry_payload_pc;
  wire       [337:0]  _zz_io_commit_0_entry_payload_uop_robPtr;
  wire       [276:0]  _zz_io_commit_0_entry_payload_uop_decoded_pc;
  wire       [4:0]    _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1;
  wire       [3:0]    _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_isa_1;
  wire       [6:0]    _zz_io_commit_0_entry_payload_uop_decoded_archDest_idx;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1;
  wire       [6:0]    _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_idx;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1;
  wire       [6:0]    _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_idx;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1;
  wire       [2:0]    _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1;
  wire       [5:0]    _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1;
  wire       [4:0]    _zz_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid;
  wire       [3:0]    _zz_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid;
  wire       [26:0]   _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1;
  wire       [17:0]   _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump;
  wire       [4:0]    _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1;
  wire       [6:0]    _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1;
  wire       [20:0]   _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1;
  wire       [17:0]   _zz_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr;
  wire       [25:0]   _zz_io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode;
  wire       [1:0]    _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1;
  wire       [33:0]   _zz_io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken;
  wire       [29:0]   _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx;
  wire       [0:0]    numToCommit;
  wire                when_ReorderBuffer_l285;
  reg        [3:0]    nextHead;
  reg        [3:0]    nextTail;
  reg        [3:0]    nextCount;
  reg        [4:0]    _zz_nextCount;
  wire       [4:0]    _zz_when_ReorderBuffer_l321;
  wire       [4:0]    _zz_when_ReorderBuffer_l321_1;
  wire                when_ReorderBuffer_l321;
  wire       [3:0]    _zz_statuses_0_genBit;
  wire       [2:0]    _zz_3;
  wire                _zz_statuses_0_genBit_1;
  wire       [31:0]   _zz_4;
  wire                _zz_5;
  wire       [4:0]    _zz_6;
  wire       [3:0]    _zz_7;
  wire       [1:0]    _zz_8;
  wire       [4:0]    _zz_9;
  wire       [1:0]    _zz_10;
  wire                _zz_11;
  wire       [4:0]    _zz_12;
  wire       [1:0]    _zz_13;
  wire                _zz_14;
  wire       [4:0]    _zz_15;
  wire       [1:0]    _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire       [31:0]   _zz_19;
  wire       [2:0]    _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire       [1:0]    _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire       [1:0]    _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire       [4:0]    _zz_40;
  wire                _zz_41;
  wire       [7:0]    _zz_42;
  wire                _zz_43;
  wire       [4:0]    _zz_44;
  wire                _zz_45;
  wire       [4:0]    _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire       [4:0]    _zz_49;
  wire       [1:0]    _zz_50;
  wire                _zz_51;
  wire       [2:0]    _zz_52;
  wire       [3:0]    _zz_53;
  wire       [1:0]    _zz_54;
  wire       [1:0]    _zz_55;
  wire       [1:0]    _zz_56;
  wire       [2:0]    _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire       [4:0]    _zz_61;
  wire       [13:0]   _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire       [19:0]   _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire       [3:0]    _zz_70;
  wire       [1:0]    _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire       [7:0]    _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire       [31:0]   _zz_78;
  wire                _zz_79;
  wire       [5:0]    _zz_80;
  wire                _zz_81;
  wire       [5:0]    _zz_82;
  wire                _zz_83;
  wire       [5:0]    _zz_84;
  wire                _zz_85;
  wire       [5:0]    _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  reg        [3:0]    _zz_90;
  wire       [15:0]   _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire       [7:0]    _zz_95;
  wire       [31:0]   _zz_96;
  wire       [7:0]    _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire       [2:0]    _zz_when_ReorderBuffer_l375;
  wire       [7:0]    _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                when_ReorderBuffer_l375;
  wire       [7:0]    _zz_statuses_0_exceptionCode;
  wire       [2:0]    _zz_when_ReorderBuffer_l375_1;
  wire       [7:0]    _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                when_ReorderBuffer_l375_1;
  wire       [7:0]    _zz_statuses_0_exceptionCode_1;
  wire       [2:0]    _zz_when_ReorderBuffer_l375_2;
  wire       [7:0]    _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire                when_ReorderBuffer_l375_2;
  wire       [7:0]    _zz_statuses_0_exceptionCode_2;
  wire       [2:0]    _zz_when_ReorderBuffer_l375_3;
  wire       [7:0]    _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                when_ReorderBuffer_l375_3;
  wire       [7:0]    _zz_statuses_0_exceptionCode_3;
  wire       [2:0]    _zz_when_ReorderBuffer_l375_4;
  wire       [7:0]    _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire                when_ReorderBuffer_l375_4;
  wire       [7:0]    _zz_statuses_0_exceptionCode_4;
  wire       [2:0]    _zz_when_ReorderBuffer_l418;
  wire       [7:0]    _zz_152;
  wire                _zz_153;
  wire                _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_1;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_2;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_3;
  reg                 when_ReorderBuffer_l418;
  wire                when_ReorderBuffer_l412;
  wire       [2:0]    _zz_when_ReorderBuffer_l418_4;
  wire       [7:0]    _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire                _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_5;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_6;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_7;
  reg                 when_ReorderBuffer_l418_1;
  wire                when_ReorderBuffer_l412_1;
  wire       [2:0]    _zz_when_ReorderBuffer_l418_8;
  wire       [7:0]    _zz_170;
  wire                _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire                _zz_174;
  wire                _zz_175;
  wire                _zz_176;
  wire                _zz_177;
  wire                _zz_178;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_9;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_10;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_11;
  reg                 when_ReorderBuffer_l418_2;
  wire                when_ReorderBuffer_l412_2;
  wire       [2:0]    _zz_when_ReorderBuffer_l418_12;
  wire       [7:0]    _zz_179;
  wire                _zz_180;
  wire                _zz_181;
  wire                _zz_182;
  wire                _zz_183;
  wire                _zz_184;
  wire                _zz_185;
  wire                _zz_186;
  wire                _zz_187;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_13;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_14;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_15;
  reg                 when_ReorderBuffer_l418_3;
  wire                when_ReorderBuffer_l412_3;
  wire       [2:0]    _zz_when_ReorderBuffer_l418_16;
  wire       [7:0]    _zz_188;
  wire                _zz_189;
  wire                _zz_190;
  wire                _zz_191;
  wire                _zz_192;
  wire                _zz_193;
  wire                _zz_194;
  wire                _zz_195;
  wire                _zz_196;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_17;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_18;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_19;
  reg                 when_ReorderBuffer_l418_4;
  wire                when_ReorderBuffer_l412_4;
  wire       [2:0]    _zz_when_ReorderBuffer_l418_20;
  wire       [7:0]    _zz_197;
  wire                _zz_198;
  wire                _zz_199;
  wire                _zz_200;
  wire                _zz_201;
  wire                _zz_202;
  wire                _zz_203;
  wire                _zz_204;
  wire                _zz_205;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_21;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_22;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_23;
  reg                 when_ReorderBuffer_l418_5;
  wire                when_ReorderBuffer_l412_5;
  wire       [2:0]    _zz_when_ReorderBuffer_l418_24;
  wire       [7:0]    _zz_206;
  wire                _zz_207;
  wire                _zz_208;
  wire                _zz_209;
  wire                _zz_210;
  wire                _zz_211;
  wire                _zz_212;
  wire                _zz_213;
  wire                _zz_214;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_25;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_26;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_27;
  reg                 when_ReorderBuffer_l418_6;
  wire                when_ReorderBuffer_l412_6;
  wire       [2:0]    _zz_when_ReorderBuffer_l418_28;
  wire       [7:0]    _zz_215;
  wire                _zz_216;
  wire                _zz_217;
  wire                _zz_218;
  wire                _zz_219;
  wire                _zz_220;
  wire                _zz_221;
  wire                _zz_222;
  wire                _zz_223;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_29;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_30;
  wire       [4:0]    _zz_when_ReorderBuffer_l418_31;
  reg                 when_ReorderBuffer_l418_7;
  wire                when_ReorderBuffer_l412_7;
  `ifndef SYNTHESIS
  reg [87:0] io_allocate_0_uopIn_decoded_uopCode_string;
  reg [151:0] io_allocate_0_uopIn_decoded_exeUnit_string;
  reg [71:0] io_allocate_0_uopIn_decoded_isa_string;
  reg [39:0] io_allocate_0_uopIn_decoded_archDest_rtype_string;
  reg [39:0] io_allocate_0_uopIn_decoded_archSrc1_rtype_string;
  reg [39:0] io_allocate_0_uopIn_decoded_archSrc2_rtype_string;
  reg [103:0] io_allocate_0_uopIn_decoded_immUsage_string;
  reg [39:0] io_allocate_0_uopIn_decoded_aluCtrl_logicOp_string;
  reg [7:0] io_allocate_0_uopIn_decoded_memCtrl_size_string;
  reg [87:0] io_allocate_0_uopIn_decoded_branchCtrl_condition_string;
  reg [39:0] io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_allocate_0_uopIn_decoded_decodeExceptionCode_string;
  reg [87:0] io_commit_0_entry_payload_uop_decoded_uopCode_string;
  reg [151:0] io_commit_0_entry_payload_uop_decoded_exeUnit_string;
  reg [71:0] io_commit_0_entry_payload_uop_decoded_isa_string;
  reg [39:0] io_commit_0_entry_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] io_commit_0_entry_payload_uop_decoded_immUsage_string;
  reg [39:0] io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] io_commit_0_entry_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string;
  reg [151:0] io_flush_payload_reason_string;
  reg [87:0] _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string;
  reg [151:0] _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string;
  reg [71:0] _zz_io_commit_0_entry_payload_uop_decoded_isa_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string;
  reg [103:0] _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string;
  reg [7:0] _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_string;
  reg [87:0] _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string;
  reg [7:0] _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string;
  reg [7:0] _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string;
  reg [7:0] _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string;
  reg [95:0] _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string;
  reg [87:0] _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string;
  reg [151:0] _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string;
  reg [71:0] _zz_io_commit_0_entry_payload_uop_decoded_isa_1_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1_string;
  reg [103:0] _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1_string;
  reg [7:0] _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1_string;
  reg [87:0] _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string;
  reg [39:0] _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1_string;
  reg [7:0] _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1_string;
  reg [7:0] _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1_string;
  reg [7:0] _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1_string;
  reg [95:0] _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1_string;
  reg [87:0] _zz_6_string;
  reg [151:0] _zz_7_string;
  reg [71:0] _zz_8_string;
  reg [39:0] _zz_10_string;
  reg [39:0] _zz_13_string;
  reg [39:0] _zz_16_string;
  reg [103:0] _zz_20_string;
  reg [39:0] _zz_25_string;
  reg [7:0] _zz_35_string;
  reg [87:0] _zz_46_string;
  reg [39:0] _zz_50_string;
  reg [7:0] _zz_54_string;
  reg [7:0] _zz_55_string;
  reg [7:0] _zz_56_string;
  reg [95:0] _zz_71_string;
  `endif

  (* ram_style = "distributed" *) reg [369:0] payloads [0:7];

  assign _zz__zz_io_allocate_0_ready = (count_reg + 4'b0000);
  assign _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx_1 = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[5 : 0];
  assign _zz_io_commit_0_entry_payload_uop_rename_physSrc2_idx = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[12 : 7];
  assign _zz_io_commit_0_entry_payload_uop_rename_physDest_idx = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[19 : 14];
  assign _zz_io_commit_0_entry_payload_uop_rename_oldPhysDest_idx = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[26 : 21];
  assign _zz_nextHead = {3'd0, numToCommit};
  assign _zz_nextTail = {3'd0, numActuallyAllocatedThisCycle};
  assign _zz_nextCount_1 = (count_reg + _zz_nextCount_2);
  assign _zz_nextCount_2 = {3'd0, numActuallyAllocatedThisCycle};
  assign _zz_nextCount_3 = {3'd0, numToCommit};
  assign _zz__zz_nextCount = (_zz_when_ReorderBuffer_l321_1 - _zz_when_ReorderBuffer_l321);
  assign _zz__zz_nextCount_1 = ({4'd0,1'b1} <<< 3'd4);
  assign _zz__zz_when_ReorderBuffer_l418_3 = {_zz__zz_when_ReorderBuffer_l418_3_1,_zz_when_ReorderBuffer_l418};
  assign _zz__zz_when_ReorderBuffer_l418_7 = {_zz__zz_when_ReorderBuffer_l418_7_1,_zz_when_ReorderBuffer_l418_4};
  assign _zz__zz_when_ReorderBuffer_l418_11 = {_zz__zz_when_ReorderBuffer_l418_11_1,_zz_when_ReorderBuffer_l418_8};
  assign _zz__zz_when_ReorderBuffer_l418_15 = {_zz__zz_when_ReorderBuffer_l418_15_1,_zz_when_ReorderBuffer_l418_12};
  assign _zz__zz_when_ReorderBuffer_l418_19 = {_zz__zz_when_ReorderBuffer_l418_19_1,_zz_when_ReorderBuffer_l418_16};
  assign _zz__zz_when_ReorderBuffer_l418_23 = {_zz__zz_when_ReorderBuffer_l418_23_1,_zz_when_ReorderBuffer_l418_20};
  assign _zz__zz_when_ReorderBuffer_l418_27 = {_zz__zz_when_ReorderBuffer_l418_27_1,_zz_when_ReorderBuffer_l418_24};
  assign _zz__zz_when_ReorderBuffer_l418_31 = {_zz__zz_when_ReorderBuffer_l418_31_1,_zz_when_ReorderBuffer_l418_28};
  assign _zz_payloads_port = {_zz_96,{_zz_95,{_zz_94,{_zz_93,{_zz_92,{_zz_91,{_zz_90,{{_zz_89,{_zz_88,{_zz_87,{_zz_86,{_zz_85,{_zz_84,{_zz_83,{_zz_82,{_zz_81,_zz_80}}}}}}}}},{{_zz_79,{_zz_78,_zz_77}},{_zz_76,{_zz_75,{_zz_74,{_zz_73,{_zz_72,{_zz_71,{{_zz_70,{_zz_69,{_zz_68,_zz_67}}},{{_zz_66,{_zz_65,{_zz_64,{_zz_63,_zz_62}}}},{{_zz_61,{_zz_60,{_zz_59,{_zz_58,{_zz_57,{_zz_56,{_zz_55,{_zz_54,_zz_53}}}}}}}},{{_zz_52,{_zz_51,{{_zz_50,_zz_49},{_zz_48,{_zz_47,_zz_46}}}}},{{_zz_45,{_zz_44,{_zz_43,{_zz_42,{_zz_41,{_zz_40,{_zz_39,{_zz_38,{_zz_37,{_zz_36,_zz_35}}}}}}}}}},{{_zz_34,{_zz_33,{_zz_32,_zz_31}}},{{_zz_30,{_zz_29,{_zz_28,{_zz_27,_zz_26}}}},{{_zz_25,{_zz_24,{_zz_23,{_zz_22,_zz_21}}}},{_zz_20,{_zz_19,{_zz_18,{_zz_17,{{_zz_16,_zz_15},{_zz_14,{{_zz_13,_zz_12},{_zz_11,{{_zz_10,_zz_9},{_zz_8,{_zz_7,{_zz_6,{_zz_5,_zz_4}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}}};
  assign _zz_numActuallyAllocatedThisCycle_1 = slotWillAllocate_0;
  assign _zz_numToCommit_1 = actualCommittedMask_0;
  assign payloads_spinal_port0 = payloads[_zz_io_commit_0_entry_status_busy];
  always @(posedge clk) begin
    if(_zz_1) begin
      payloads[_zz_3] <= _zz_payloads_port;
    end
  end

  always @(*) begin
    case(_zz_numActuallyAllocatedThisCycle_1)
      1'b0 : _zz_numActuallyAllocatedThisCycle = 1'b0;
      default : _zz_numActuallyAllocatedThisCycle = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_io_commit_0_entry_status_busy)
      3'b000 : begin
        _zz__zz_io_commit_0_entry_status_done = statuses_0_done;
        _zz__zz_io_commit_0_entry_status_genBit = statuses_0_genBit;
        _zz_io_commit_0_entry_status_busy_1 = statuses_0_busy;
        _zz_io_commit_0_entry_status_isMispredictedBranch = statuses_0_isMispredictedBranch;
        _zz_io_commit_0_entry_status_isTaken = statuses_0_isTaken;
        _zz_io_commit_0_entry_status_result = statuses_0_result;
        _zz_io_commit_0_entry_status_hasException = statuses_0_hasException;
        _zz_io_commit_0_entry_status_exceptionCode = statuses_0_exceptionCode;
      end
      3'b001 : begin
        _zz__zz_io_commit_0_entry_status_done = statuses_1_done;
        _zz__zz_io_commit_0_entry_status_genBit = statuses_1_genBit;
        _zz_io_commit_0_entry_status_busy_1 = statuses_1_busy;
        _zz_io_commit_0_entry_status_isMispredictedBranch = statuses_1_isMispredictedBranch;
        _zz_io_commit_0_entry_status_isTaken = statuses_1_isTaken;
        _zz_io_commit_0_entry_status_result = statuses_1_result;
        _zz_io_commit_0_entry_status_hasException = statuses_1_hasException;
        _zz_io_commit_0_entry_status_exceptionCode = statuses_1_exceptionCode;
      end
      3'b010 : begin
        _zz__zz_io_commit_0_entry_status_done = statuses_2_done;
        _zz__zz_io_commit_0_entry_status_genBit = statuses_2_genBit;
        _zz_io_commit_0_entry_status_busy_1 = statuses_2_busy;
        _zz_io_commit_0_entry_status_isMispredictedBranch = statuses_2_isMispredictedBranch;
        _zz_io_commit_0_entry_status_isTaken = statuses_2_isTaken;
        _zz_io_commit_0_entry_status_result = statuses_2_result;
        _zz_io_commit_0_entry_status_hasException = statuses_2_hasException;
        _zz_io_commit_0_entry_status_exceptionCode = statuses_2_exceptionCode;
      end
      3'b011 : begin
        _zz__zz_io_commit_0_entry_status_done = statuses_3_done;
        _zz__zz_io_commit_0_entry_status_genBit = statuses_3_genBit;
        _zz_io_commit_0_entry_status_busy_1 = statuses_3_busy;
        _zz_io_commit_0_entry_status_isMispredictedBranch = statuses_3_isMispredictedBranch;
        _zz_io_commit_0_entry_status_isTaken = statuses_3_isTaken;
        _zz_io_commit_0_entry_status_result = statuses_3_result;
        _zz_io_commit_0_entry_status_hasException = statuses_3_hasException;
        _zz_io_commit_0_entry_status_exceptionCode = statuses_3_exceptionCode;
      end
      3'b100 : begin
        _zz__zz_io_commit_0_entry_status_done = statuses_4_done;
        _zz__zz_io_commit_0_entry_status_genBit = statuses_4_genBit;
        _zz_io_commit_0_entry_status_busy_1 = statuses_4_busy;
        _zz_io_commit_0_entry_status_isMispredictedBranch = statuses_4_isMispredictedBranch;
        _zz_io_commit_0_entry_status_isTaken = statuses_4_isTaken;
        _zz_io_commit_0_entry_status_result = statuses_4_result;
        _zz_io_commit_0_entry_status_hasException = statuses_4_hasException;
        _zz_io_commit_0_entry_status_exceptionCode = statuses_4_exceptionCode;
      end
      3'b101 : begin
        _zz__zz_io_commit_0_entry_status_done = statuses_5_done;
        _zz__zz_io_commit_0_entry_status_genBit = statuses_5_genBit;
        _zz_io_commit_0_entry_status_busy_1 = statuses_5_busy;
        _zz_io_commit_0_entry_status_isMispredictedBranch = statuses_5_isMispredictedBranch;
        _zz_io_commit_0_entry_status_isTaken = statuses_5_isTaken;
        _zz_io_commit_0_entry_status_result = statuses_5_result;
        _zz_io_commit_0_entry_status_hasException = statuses_5_hasException;
        _zz_io_commit_0_entry_status_exceptionCode = statuses_5_exceptionCode;
      end
      3'b110 : begin
        _zz__zz_io_commit_0_entry_status_done = statuses_6_done;
        _zz__zz_io_commit_0_entry_status_genBit = statuses_6_genBit;
        _zz_io_commit_0_entry_status_busy_1 = statuses_6_busy;
        _zz_io_commit_0_entry_status_isMispredictedBranch = statuses_6_isMispredictedBranch;
        _zz_io_commit_0_entry_status_isTaken = statuses_6_isTaken;
        _zz_io_commit_0_entry_status_result = statuses_6_result;
        _zz_io_commit_0_entry_status_hasException = statuses_6_hasException;
        _zz_io_commit_0_entry_status_exceptionCode = statuses_6_exceptionCode;
      end
      default : begin
        _zz__zz_io_commit_0_entry_status_done = statuses_7_done;
        _zz__zz_io_commit_0_entry_status_genBit = statuses_7_genBit;
        _zz_io_commit_0_entry_status_busy_1 = statuses_7_busy;
        _zz_io_commit_0_entry_status_isMispredictedBranch = statuses_7_isMispredictedBranch;
        _zz_io_commit_0_entry_status_isTaken = statuses_7_isTaken;
        _zz_io_commit_0_entry_status_result = statuses_7_result;
        _zz_io_commit_0_entry_status_hasException = statuses_7_hasException;
        _zz_io_commit_0_entry_status_exceptionCode = statuses_7_exceptionCode;
      end
    endcase
  end

  always @(*) begin
    case(_zz_numToCommit_1)
      1'b0 : _zz_numToCommit = 1'b0;
      default : _zz_numToCommit = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l375)
      3'b000 : begin
        _zz_when_ReorderBuffer_l375_5 = statuses_0_genBit;
        _zz__zz_statuses_0_exceptionCode = statuses_0_exceptionCode;
      end
      3'b001 : begin
        _zz_when_ReorderBuffer_l375_5 = statuses_1_genBit;
        _zz__zz_statuses_0_exceptionCode = statuses_1_exceptionCode;
      end
      3'b010 : begin
        _zz_when_ReorderBuffer_l375_5 = statuses_2_genBit;
        _zz__zz_statuses_0_exceptionCode = statuses_2_exceptionCode;
      end
      3'b011 : begin
        _zz_when_ReorderBuffer_l375_5 = statuses_3_genBit;
        _zz__zz_statuses_0_exceptionCode = statuses_3_exceptionCode;
      end
      3'b100 : begin
        _zz_when_ReorderBuffer_l375_5 = statuses_4_genBit;
        _zz__zz_statuses_0_exceptionCode = statuses_4_exceptionCode;
      end
      3'b101 : begin
        _zz_when_ReorderBuffer_l375_5 = statuses_5_genBit;
        _zz__zz_statuses_0_exceptionCode = statuses_5_exceptionCode;
      end
      3'b110 : begin
        _zz_when_ReorderBuffer_l375_5 = statuses_6_genBit;
        _zz__zz_statuses_0_exceptionCode = statuses_6_exceptionCode;
      end
      default : begin
        _zz_when_ReorderBuffer_l375_5 = statuses_7_genBit;
        _zz__zz_statuses_0_exceptionCode = statuses_7_exceptionCode;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l375_1)
      3'b000 : begin
        _zz_when_ReorderBuffer_l375_1_1 = statuses_0_genBit;
        _zz__zz_statuses_0_exceptionCode_1 = statuses_0_exceptionCode;
      end
      3'b001 : begin
        _zz_when_ReorderBuffer_l375_1_1 = statuses_1_genBit;
        _zz__zz_statuses_0_exceptionCode_1 = statuses_1_exceptionCode;
      end
      3'b010 : begin
        _zz_when_ReorderBuffer_l375_1_1 = statuses_2_genBit;
        _zz__zz_statuses_0_exceptionCode_1 = statuses_2_exceptionCode;
      end
      3'b011 : begin
        _zz_when_ReorderBuffer_l375_1_1 = statuses_3_genBit;
        _zz__zz_statuses_0_exceptionCode_1 = statuses_3_exceptionCode;
      end
      3'b100 : begin
        _zz_when_ReorderBuffer_l375_1_1 = statuses_4_genBit;
        _zz__zz_statuses_0_exceptionCode_1 = statuses_4_exceptionCode;
      end
      3'b101 : begin
        _zz_when_ReorderBuffer_l375_1_1 = statuses_5_genBit;
        _zz__zz_statuses_0_exceptionCode_1 = statuses_5_exceptionCode;
      end
      3'b110 : begin
        _zz_when_ReorderBuffer_l375_1_1 = statuses_6_genBit;
        _zz__zz_statuses_0_exceptionCode_1 = statuses_6_exceptionCode;
      end
      default : begin
        _zz_when_ReorderBuffer_l375_1_1 = statuses_7_genBit;
        _zz__zz_statuses_0_exceptionCode_1 = statuses_7_exceptionCode;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l375_2)
      3'b000 : begin
        _zz_when_ReorderBuffer_l375_2_1 = statuses_0_genBit;
        _zz__zz_statuses_0_exceptionCode_2 = statuses_0_exceptionCode;
      end
      3'b001 : begin
        _zz_when_ReorderBuffer_l375_2_1 = statuses_1_genBit;
        _zz__zz_statuses_0_exceptionCode_2 = statuses_1_exceptionCode;
      end
      3'b010 : begin
        _zz_when_ReorderBuffer_l375_2_1 = statuses_2_genBit;
        _zz__zz_statuses_0_exceptionCode_2 = statuses_2_exceptionCode;
      end
      3'b011 : begin
        _zz_when_ReorderBuffer_l375_2_1 = statuses_3_genBit;
        _zz__zz_statuses_0_exceptionCode_2 = statuses_3_exceptionCode;
      end
      3'b100 : begin
        _zz_when_ReorderBuffer_l375_2_1 = statuses_4_genBit;
        _zz__zz_statuses_0_exceptionCode_2 = statuses_4_exceptionCode;
      end
      3'b101 : begin
        _zz_when_ReorderBuffer_l375_2_1 = statuses_5_genBit;
        _zz__zz_statuses_0_exceptionCode_2 = statuses_5_exceptionCode;
      end
      3'b110 : begin
        _zz_when_ReorderBuffer_l375_2_1 = statuses_6_genBit;
        _zz__zz_statuses_0_exceptionCode_2 = statuses_6_exceptionCode;
      end
      default : begin
        _zz_when_ReorderBuffer_l375_2_1 = statuses_7_genBit;
        _zz__zz_statuses_0_exceptionCode_2 = statuses_7_exceptionCode;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l375_3)
      3'b000 : begin
        _zz_when_ReorderBuffer_l375_3_1 = statuses_0_genBit;
        _zz__zz_statuses_0_exceptionCode_3 = statuses_0_exceptionCode;
      end
      3'b001 : begin
        _zz_when_ReorderBuffer_l375_3_1 = statuses_1_genBit;
        _zz__zz_statuses_0_exceptionCode_3 = statuses_1_exceptionCode;
      end
      3'b010 : begin
        _zz_when_ReorderBuffer_l375_3_1 = statuses_2_genBit;
        _zz__zz_statuses_0_exceptionCode_3 = statuses_2_exceptionCode;
      end
      3'b011 : begin
        _zz_when_ReorderBuffer_l375_3_1 = statuses_3_genBit;
        _zz__zz_statuses_0_exceptionCode_3 = statuses_3_exceptionCode;
      end
      3'b100 : begin
        _zz_when_ReorderBuffer_l375_3_1 = statuses_4_genBit;
        _zz__zz_statuses_0_exceptionCode_3 = statuses_4_exceptionCode;
      end
      3'b101 : begin
        _zz_when_ReorderBuffer_l375_3_1 = statuses_5_genBit;
        _zz__zz_statuses_0_exceptionCode_3 = statuses_5_exceptionCode;
      end
      3'b110 : begin
        _zz_when_ReorderBuffer_l375_3_1 = statuses_6_genBit;
        _zz__zz_statuses_0_exceptionCode_3 = statuses_6_exceptionCode;
      end
      default : begin
        _zz_when_ReorderBuffer_l375_3_1 = statuses_7_genBit;
        _zz__zz_statuses_0_exceptionCode_3 = statuses_7_exceptionCode;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l375_4)
      3'b000 : begin
        _zz_when_ReorderBuffer_l375_4_1 = statuses_0_genBit;
        _zz__zz_statuses_0_exceptionCode_4 = statuses_0_exceptionCode;
      end
      3'b001 : begin
        _zz_when_ReorderBuffer_l375_4_1 = statuses_1_genBit;
        _zz__zz_statuses_0_exceptionCode_4 = statuses_1_exceptionCode;
      end
      3'b010 : begin
        _zz_when_ReorderBuffer_l375_4_1 = statuses_2_genBit;
        _zz__zz_statuses_0_exceptionCode_4 = statuses_2_exceptionCode;
      end
      3'b011 : begin
        _zz_when_ReorderBuffer_l375_4_1 = statuses_3_genBit;
        _zz__zz_statuses_0_exceptionCode_4 = statuses_3_exceptionCode;
      end
      3'b100 : begin
        _zz_when_ReorderBuffer_l375_4_1 = statuses_4_genBit;
        _zz__zz_statuses_0_exceptionCode_4 = statuses_4_exceptionCode;
      end
      3'b101 : begin
        _zz_when_ReorderBuffer_l375_4_1 = statuses_5_genBit;
        _zz__zz_statuses_0_exceptionCode_4 = statuses_5_exceptionCode;
      end
      3'b110 : begin
        _zz_when_ReorderBuffer_l375_4_1 = statuses_6_genBit;
        _zz__zz_statuses_0_exceptionCode_4 = statuses_6_exceptionCode;
      end
      default : begin
        _zz_when_ReorderBuffer_l375_4_1 = statuses_7_genBit;
        _zz__zz_statuses_0_exceptionCode_4 = statuses_7_exceptionCode;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l418)
      3'b000 : _zz__zz_when_ReorderBuffer_l418_3_1 = statuses_0_genBit;
      3'b001 : _zz__zz_when_ReorderBuffer_l418_3_1 = statuses_1_genBit;
      3'b010 : _zz__zz_when_ReorderBuffer_l418_3_1 = statuses_2_genBit;
      3'b011 : _zz__zz_when_ReorderBuffer_l418_3_1 = statuses_3_genBit;
      3'b100 : _zz__zz_when_ReorderBuffer_l418_3_1 = statuses_4_genBit;
      3'b101 : _zz__zz_when_ReorderBuffer_l418_3_1 = statuses_5_genBit;
      3'b110 : _zz__zz_when_ReorderBuffer_l418_3_1 = statuses_6_genBit;
      default : _zz__zz_when_ReorderBuffer_l418_3_1 = statuses_7_genBit;
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l418_4)
      3'b000 : _zz__zz_when_ReorderBuffer_l418_7_1 = statuses_0_genBit;
      3'b001 : _zz__zz_when_ReorderBuffer_l418_7_1 = statuses_1_genBit;
      3'b010 : _zz__zz_when_ReorderBuffer_l418_7_1 = statuses_2_genBit;
      3'b011 : _zz__zz_when_ReorderBuffer_l418_7_1 = statuses_3_genBit;
      3'b100 : _zz__zz_when_ReorderBuffer_l418_7_1 = statuses_4_genBit;
      3'b101 : _zz__zz_when_ReorderBuffer_l418_7_1 = statuses_5_genBit;
      3'b110 : _zz__zz_when_ReorderBuffer_l418_7_1 = statuses_6_genBit;
      default : _zz__zz_when_ReorderBuffer_l418_7_1 = statuses_7_genBit;
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l418_8)
      3'b000 : _zz__zz_when_ReorderBuffer_l418_11_1 = statuses_0_genBit;
      3'b001 : _zz__zz_when_ReorderBuffer_l418_11_1 = statuses_1_genBit;
      3'b010 : _zz__zz_when_ReorderBuffer_l418_11_1 = statuses_2_genBit;
      3'b011 : _zz__zz_when_ReorderBuffer_l418_11_1 = statuses_3_genBit;
      3'b100 : _zz__zz_when_ReorderBuffer_l418_11_1 = statuses_4_genBit;
      3'b101 : _zz__zz_when_ReorderBuffer_l418_11_1 = statuses_5_genBit;
      3'b110 : _zz__zz_when_ReorderBuffer_l418_11_1 = statuses_6_genBit;
      default : _zz__zz_when_ReorderBuffer_l418_11_1 = statuses_7_genBit;
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l418_12)
      3'b000 : _zz__zz_when_ReorderBuffer_l418_15_1 = statuses_0_genBit;
      3'b001 : _zz__zz_when_ReorderBuffer_l418_15_1 = statuses_1_genBit;
      3'b010 : _zz__zz_when_ReorderBuffer_l418_15_1 = statuses_2_genBit;
      3'b011 : _zz__zz_when_ReorderBuffer_l418_15_1 = statuses_3_genBit;
      3'b100 : _zz__zz_when_ReorderBuffer_l418_15_1 = statuses_4_genBit;
      3'b101 : _zz__zz_when_ReorderBuffer_l418_15_1 = statuses_5_genBit;
      3'b110 : _zz__zz_when_ReorderBuffer_l418_15_1 = statuses_6_genBit;
      default : _zz__zz_when_ReorderBuffer_l418_15_1 = statuses_7_genBit;
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l418_16)
      3'b000 : _zz__zz_when_ReorderBuffer_l418_19_1 = statuses_0_genBit;
      3'b001 : _zz__zz_when_ReorderBuffer_l418_19_1 = statuses_1_genBit;
      3'b010 : _zz__zz_when_ReorderBuffer_l418_19_1 = statuses_2_genBit;
      3'b011 : _zz__zz_when_ReorderBuffer_l418_19_1 = statuses_3_genBit;
      3'b100 : _zz__zz_when_ReorderBuffer_l418_19_1 = statuses_4_genBit;
      3'b101 : _zz__zz_when_ReorderBuffer_l418_19_1 = statuses_5_genBit;
      3'b110 : _zz__zz_when_ReorderBuffer_l418_19_1 = statuses_6_genBit;
      default : _zz__zz_when_ReorderBuffer_l418_19_1 = statuses_7_genBit;
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l418_20)
      3'b000 : _zz__zz_when_ReorderBuffer_l418_23_1 = statuses_0_genBit;
      3'b001 : _zz__zz_when_ReorderBuffer_l418_23_1 = statuses_1_genBit;
      3'b010 : _zz__zz_when_ReorderBuffer_l418_23_1 = statuses_2_genBit;
      3'b011 : _zz__zz_when_ReorderBuffer_l418_23_1 = statuses_3_genBit;
      3'b100 : _zz__zz_when_ReorderBuffer_l418_23_1 = statuses_4_genBit;
      3'b101 : _zz__zz_when_ReorderBuffer_l418_23_1 = statuses_5_genBit;
      3'b110 : _zz__zz_when_ReorderBuffer_l418_23_1 = statuses_6_genBit;
      default : _zz__zz_when_ReorderBuffer_l418_23_1 = statuses_7_genBit;
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l418_24)
      3'b000 : _zz__zz_when_ReorderBuffer_l418_27_1 = statuses_0_genBit;
      3'b001 : _zz__zz_when_ReorderBuffer_l418_27_1 = statuses_1_genBit;
      3'b010 : _zz__zz_when_ReorderBuffer_l418_27_1 = statuses_2_genBit;
      3'b011 : _zz__zz_when_ReorderBuffer_l418_27_1 = statuses_3_genBit;
      3'b100 : _zz__zz_when_ReorderBuffer_l418_27_1 = statuses_4_genBit;
      3'b101 : _zz__zz_when_ReorderBuffer_l418_27_1 = statuses_5_genBit;
      3'b110 : _zz__zz_when_ReorderBuffer_l418_27_1 = statuses_6_genBit;
      default : _zz__zz_when_ReorderBuffer_l418_27_1 = statuses_7_genBit;
    endcase
  end

  always @(*) begin
    case(_zz_when_ReorderBuffer_l418_28)
      3'b000 : _zz__zz_when_ReorderBuffer_l418_31_1 = statuses_0_genBit;
      3'b001 : _zz__zz_when_ReorderBuffer_l418_31_1 = statuses_1_genBit;
      3'b010 : _zz__zz_when_ReorderBuffer_l418_31_1 = statuses_2_genBit;
      3'b011 : _zz__zz_when_ReorderBuffer_l418_31_1 = statuses_3_genBit;
      3'b100 : _zz__zz_when_ReorderBuffer_l418_31_1 = statuses_4_genBit;
      3'b101 : _zz__zz_when_ReorderBuffer_l418_31_1 = statuses_5_genBit;
      3'b110 : _zz__zz_when_ReorderBuffer_l418_31_1 = statuses_6_genBit;
      default : _zz__zz_when_ReorderBuffer_l418_31_1 = statuses_7_genBit;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_uopCode)
      BaseUopCode_NOP : io_allocate_0_uopIn_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_allocate_0_uopIn_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_allocate_0_uopIn_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_allocate_0_uopIn_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_allocate_0_uopIn_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_allocate_0_uopIn_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_allocate_0_uopIn_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_allocate_0_uopIn_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_allocate_0_uopIn_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_allocate_0_uopIn_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_allocate_0_uopIn_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_allocate_0_uopIn_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_allocate_0_uopIn_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_allocate_0_uopIn_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_allocate_0_uopIn_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_allocate_0_uopIn_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_allocate_0_uopIn_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_allocate_0_uopIn_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_allocate_0_uopIn_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_allocate_0_uopIn_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_allocate_0_uopIn_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_allocate_0_uopIn_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_allocate_0_uopIn_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_allocate_0_uopIn_decoded_uopCode_string = "IDLE       ";
      default : io_allocate_0_uopIn_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_exeUnit)
      ExeUnitType_NONE : io_allocate_0_uopIn_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_allocate_0_uopIn_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_allocate_0_uopIn_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_allocate_0_uopIn_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_allocate_0_uopIn_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_allocate_0_uopIn_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_allocate_0_uopIn_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_allocate_0_uopIn_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_allocate_0_uopIn_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_allocate_0_uopIn_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_isa)
      IsaType_UNKNOWN : io_allocate_0_uopIn_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_allocate_0_uopIn_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : io_allocate_0_uopIn_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_allocate_0_uopIn_decoded_isa_string = "LOONGARCH";
      default : io_allocate_0_uopIn_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_archDest_rtype)
      ArchRegType_GPR : io_allocate_0_uopIn_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocate_0_uopIn_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocate_0_uopIn_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocate_0_uopIn_decoded_archDest_rtype_string = "LA_CF";
      default : io_allocate_0_uopIn_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_archSrc1_rtype)
      ArchRegType_GPR : io_allocate_0_uopIn_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocate_0_uopIn_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocate_0_uopIn_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocate_0_uopIn_decoded_archSrc1_rtype_string = "LA_CF";
      default : io_allocate_0_uopIn_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_archSrc2_rtype)
      ArchRegType_GPR : io_allocate_0_uopIn_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocate_0_uopIn_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocate_0_uopIn_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocate_0_uopIn_decoded_archSrc2_rtype_string = "LA_CF";
      default : io_allocate_0_uopIn_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_immUsage)
      ImmUsageType_NONE : io_allocate_0_uopIn_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_allocate_0_uopIn_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_allocate_0_uopIn_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_allocate_0_uopIn_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_allocate_0_uopIn_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_allocate_0_uopIn_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_allocate_0_uopIn_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : io_allocate_0_uopIn_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_aluCtrl_logicOp)
      LogicOp_NONE : io_allocate_0_uopIn_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_allocate_0_uopIn_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_allocate_0_uopIn_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_allocate_0_uopIn_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : io_allocate_0_uopIn_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_memCtrl_size)
      MemAccessSize_B : io_allocate_0_uopIn_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : io_allocate_0_uopIn_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : io_allocate_0_uopIn_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : io_allocate_0_uopIn_decoded_memCtrl_size_string = "D";
      default : io_allocate_0_uopIn_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_branchCtrl_condition)
      BranchCondition_NUL : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_allocate_0_uopIn_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_allocate_0_uopIn_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : io_allocate_0_uopIn_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_allocate_0_uopIn_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_allocate_0_uopIn_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_allocate_0_uopIn_decoded_decodeExceptionCode_string = "OK          ";
      default : io_allocate_0_uopIn_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : io_commit_0_entry_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : io_commit_0_entry_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : io_commit_0_entry_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : io_commit_0_entry_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : io_commit_0_entry_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : io_commit_0_entry_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : io_commit_0_entry_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : io_commit_0_entry_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : io_commit_0_entry_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : io_commit_0_entry_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : io_commit_0_entry_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : io_commit_0_entry_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : io_commit_0_entry_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : io_commit_0_entry_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : io_commit_0_entry_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : io_commit_0_entry_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : io_commit_0_entry_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : io_commit_0_entry_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : io_commit_0_entry_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : io_commit_0_entry_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : io_commit_0_entry_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : io_commit_0_entry_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : io_commit_0_entry_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : io_commit_0_entry_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : io_commit_0_entry_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : io_commit_0_entry_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_isa)
      IsaType_UNKNOWN : io_commit_0_entry_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : io_commit_0_entry_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : io_commit_0_entry_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : io_commit_0_entry_payload_uop_decoded_isa_string = "LOONGARCH";
      default : io_commit_0_entry_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : io_commit_0_entry_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_commit_0_entry_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_commit_0_entry_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_commit_0_entry_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_commit_0_entry_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_commit_0_entry_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_commit_0_entry_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : io_commit_0_entry_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "D";
      default : io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(io_commit_0_entry_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_flush_payload_reason)
      FlushReason_NONE : io_flush_payload_reason_string = "NONE               ";
      FlushReason_FULL_FLUSH : io_flush_payload_reason_string = "FULL_FLUSH         ";
      FlushReason_ROLLBACK_TO_ROB_IDX : io_flush_payload_reason_string = "ROLLBACK_TO_ROB_IDX";
      default : io_flush_payload_reason_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_uopCode)
      BaseUopCode_NOP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "NOP        ";
      BaseUopCode_ILLEGAL : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "ILLEGAL    ";
      BaseUopCode_ALU : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "ALU        ";
      BaseUopCode_SHIFT : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "SHIFT      ";
      BaseUopCode_MUL : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "MUL        ";
      BaseUopCode_DIV : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "DIV        ";
      BaseUopCode_LOAD : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "LOAD       ";
      BaseUopCode_STORE : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "STORE      ";
      BaseUopCode_ATOMIC : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "PREFETCH   ";
      BaseUopCode_BRANCH : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "LA_TLB     ";
      BaseUopCode_IDLE : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "IDLE       ";
      default : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_exeUnit)
      ExeUnitType_NONE : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "NONE               ";
      ExeUnitType_ALU_INT : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "DIV_INT            ";
      ExeUnitType_MEM : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "MEM                ";
      ExeUnitType_BRU : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "BRU                ";
      ExeUnitType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "FPU_DIV_SQRT       ";
      default : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_isa)
      IsaType_UNKNOWN : _zz_io_commit_0_entry_payload_uop_decoded_isa_string = "UNKNOWN  ";
      IsaType_DEMO : _zz_io_commit_0_entry_payload_uop_decoded_isa_string = "DEMO     ";
      IsaType_RISCV : _zz_io_commit_0_entry_payload_uop_decoded_isa_string = "RISCV    ";
      IsaType_LOONGARCH : _zz_io_commit_0_entry_payload_uop_decoded_isa_string = "LOONGARCH";
      default : _zz_io_commit_0_entry_payload_uop_decoded_isa_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype)
      ArchRegType_GPR : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "LA_CF";
      default : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype)
      ArchRegType_GPR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "LA_CF";
      default : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype)
      ArchRegType_GPR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "LA_CF";
      default : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_immUsage)
      ImmUsageType_NONE : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string = "JUMP_OFFSET  ";
      default : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp)
      LogicOp_NONE : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "XOR_1";
      default : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size)
      MemAccessSize_B : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "B";
      MemAccessSize_H : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "H";
      MemAccessSize_W : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "W";
      MemAccessSize_D : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "D";
      default : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition)
      BranchCondition_NUL : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "NUL        ";
      BranchCondition_EQ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "EQ         ";
      BranchCondition_NE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "NE         ";
      BranchCondition_LT : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LT         ";
      BranchCondition_GE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "GE         ";
      BranchCondition_LTU : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LTU        ";
      BranchCondition_GEU : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "GEU        ";
      BranchCondition_EQZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "EQZ        ";
      BranchCondition_NEZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "NEZ        ";
      BranchCondition_LTZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LTZ        ";
      BranchCondition_GEZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "GEZ        ";
      BranchCondition_GTZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "GTZ        ";
      BranchCondition_LEZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_NE       ";
      BranchCondition_F_LT : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_LT       ";
      BranchCondition_F_LE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_LE       ";
      BranchCondition_F_UN : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "LA_CF_FALSE";
      default : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype)
      ArchRegType_GPR : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "GPR  ";
      ArchRegType_FPR : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "FPR  ";
      ArchRegType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "LA_CF";
      default : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1)
      MemAccessSize_B : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "B";
      MemAccessSize_H : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "H";
      MemAccessSize_W : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "W";
      MemAccessSize_D : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "D";
      default : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2)
      MemAccessSize_B : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "B";
      MemAccessSize_H : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "H";
      MemAccessSize_W : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "W";
      MemAccessSize_D : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "D";
      default : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest)
      MemAccessSize_B : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "B";
      MemAccessSize_H : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "H";
      MemAccessSize_W : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "W";
      MemAccessSize_D : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "D";
      default : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode)
      DecodeExCode_INVALID : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "DECODE_ERROR";
      DecodeExCode_OK : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "OK          ";
      default : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_uopCode_1)
      BaseUopCode_NOP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "NOP        ";
      BaseUopCode_ILLEGAL : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "ILLEGAL    ";
      BaseUopCode_ALU : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "ALU        ";
      BaseUopCode_SHIFT : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "SHIFT      ";
      BaseUopCode_MUL : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "MUL        ";
      BaseUopCode_DIV : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "DIV        ";
      BaseUopCode_LOAD : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "LOAD       ";
      BaseUopCode_STORE : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "STORE      ";
      BaseUopCode_ATOMIC : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "PREFETCH   ";
      BaseUopCode_BRANCH : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "LA_TLB     ";
      BaseUopCode_IDLE : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "IDLE       ";
      default : _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1)
      ExeUnitType_NONE : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "NONE               ";
      ExeUnitType_ALU_INT : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "DIV_INT            ";
      ExeUnitType_MEM : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "MEM                ";
      ExeUnitType_BRU : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "BRU                ";
      ExeUnitType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "FPU_DIV_SQRT       ";
      default : _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_isa_1)
      IsaType_UNKNOWN : _zz_io_commit_0_entry_payload_uop_decoded_isa_1_string = "UNKNOWN  ";
      IsaType_DEMO : _zz_io_commit_0_entry_payload_uop_decoded_isa_1_string = "DEMO     ";
      IsaType_RISCV : _zz_io_commit_0_entry_payload_uop_decoded_isa_1_string = "RISCV    ";
      IsaType_LOONGARCH : _zz_io_commit_0_entry_payload_uop_decoded_isa_1_string = "LOONGARCH";
      default : _zz_io_commit_0_entry_payload_uop_decoded_isa_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1)
      ArchRegType_GPR : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1_string = "GPR  ";
      ArchRegType_FPR : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1_string = "FPR  ";
      ArchRegType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1_string = "LA_CF";
      default : _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1)
      ArchRegType_GPR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1_string = "GPR  ";
      ArchRegType_FPR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1_string = "FPR  ";
      ArchRegType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1_string = "LA_CF";
      default : _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1)
      ArchRegType_GPR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1_string = "GPR  ";
      ArchRegType_FPR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1_string = "FPR  ";
      ArchRegType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1_string = "LA_CF";
      default : _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_immUsage_1)
      ImmUsageType_NONE : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string = "JUMP_OFFSET  ";
      default : _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1)
      LogicOp_NONE : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1_string = "NONE ";
      LogicOp_AND_1 : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1_string = "AND_1";
      LogicOp_OR_1 : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1_string = "XOR_1";
      default : _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1)
      MemAccessSize_B : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1_string = "B";
      MemAccessSize_H : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1_string = "H";
      MemAccessSize_W : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1_string = "W";
      MemAccessSize_D : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1_string = "D";
      default : _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1)
      BranchCondition_NUL : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "NUL        ";
      BranchCondition_EQ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "EQ         ";
      BranchCondition_NE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "NE         ";
      BranchCondition_LT : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "LT         ";
      BranchCondition_GE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "GE         ";
      BranchCondition_LTU : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "LTU        ";
      BranchCondition_GEU : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "GEU        ";
      BranchCondition_EQZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "EQZ        ";
      BranchCondition_NEZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "NEZ        ";
      BranchCondition_LTZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "LTZ        ";
      BranchCondition_GEZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "GEZ        ";
      BranchCondition_GTZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "GTZ        ";
      BranchCondition_LEZ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "F_NE       ";
      BranchCondition_F_LT : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "F_LT       ";
      BranchCondition_F_LE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "F_LE       ";
      BranchCondition_F_UN : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "LA_CF_FALSE";
      default : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1)
      ArchRegType_GPR : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1_string = "GPR  ";
      ArchRegType_FPR : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1_string = "FPR  ";
      ArchRegType_CSR : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1_string = "CSR  ";
      ArchRegType_LA_CF : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1_string = "LA_CF";
      default : _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1)
      MemAccessSize_B : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1_string = "B";
      MemAccessSize_H : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1_string = "H";
      MemAccessSize_W : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1_string = "W";
      MemAccessSize_D : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1_string = "D";
      default : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1)
      MemAccessSize_B : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1_string = "B";
      MemAccessSize_H : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1_string = "H";
      MemAccessSize_W : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1_string = "W";
      MemAccessSize_D : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1_string = "D";
      default : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1)
      MemAccessSize_B : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1_string = "B";
      MemAccessSize_H : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1_string = "H";
      MemAccessSize_W : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1_string = "W";
      MemAccessSize_D : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1_string = "D";
      default : _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1)
      DecodeExCode_INVALID : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1_string = "DECODE_ERROR";
      DecodeExCode_OK : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1_string = "OK          ";
      default : _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_6)
      BaseUopCode_NOP : _zz_6_string = "NOP        ";
      BaseUopCode_ILLEGAL : _zz_6_string = "ILLEGAL    ";
      BaseUopCode_ALU : _zz_6_string = "ALU        ";
      BaseUopCode_SHIFT : _zz_6_string = "SHIFT      ";
      BaseUopCode_MUL : _zz_6_string = "MUL        ";
      BaseUopCode_DIV : _zz_6_string = "DIV        ";
      BaseUopCode_LOAD : _zz_6_string = "LOAD       ";
      BaseUopCode_STORE : _zz_6_string = "STORE      ";
      BaseUopCode_ATOMIC : _zz_6_string = "ATOMIC     ";
      BaseUopCode_MEM_BARRIER : _zz_6_string = "MEM_BARRIER";
      BaseUopCode_PREFETCH : _zz_6_string = "PREFETCH   ";
      BaseUopCode_BRANCH : _zz_6_string = "BRANCH     ";
      BaseUopCode_JUMP_REG : _zz_6_string = "JUMP_REG   ";
      BaseUopCode_JUMP_IMM : _zz_6_string = "JUMP_IMM   ";
      BaseUopCode_SYSTEM_OP : _zz_6_string = "SYSTEM_OP  ";
      BaseUopCode_CSR_ACCESS : _zz_6_string = "CSR_ACCESS ";
      BaseUopCode_FPU_ALU : _zz_6_string = "FPU_ALU    ";
      BaseUopCode_FPU_CVT : _zz_6_string = "FPU_CVT    ";
      BaseUopCode_FPU_CMP : _zz_6_string = "FPU_CMP    ";
      BaseUopCode_FPU_SEL : _zz_6_string = "FPU_SEL    ";
      BaseUopCode_LA_BITMANIP : _zz_6_string = "LA_BITMANIP";
      BaseUopCode_LA_CACOP : _zz_6_string = "LA_CACOP   ";
      BaseUopCode_LA_TLB : _zz_6_string = "LA_TLB     ";
      BaseUopCode_IDLE : _zz_6_string = "IDLE       ";
      default : _zz_6_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_7)
      ExeUnitType_NONE : _zz_7_string = "NONE               ";
      ExeUnitType_ALU_INT : _zz_7_string = "ALU_INT            ";
      ExeUnitType_MUL_INT : _zz_7_string = "MUL_INT            ";
      ExeUnitType_DIV_INT : _zz_7_string = "DIV_INT            ";
      ExeUnitType_MEM : _zz_7_string = "MEM                ";
      ExeUnitType_BRU : _zz_7_string = "BRU                ";
      ExeUnitType_CSR : _zz_7_string = "CSR                ";
      ExeUnitType_FPU_ADD_MUL_CVT_CMP : _zz_7_string = "FPU_ADD_MUL_CVT_CMP";
      ExeUnitType_FPU_DIV_SQRT : _zz_7_string = "FPU_DIV_SQRT       ";
      default : _zz_7_string = "???????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_8)
      IsaType_UNKNOWN : _zz_8_string = "UNKNOWN  ";
      IsaType_DEMO : _zz_8_string = "DEMO     ";
      IsaType_RISCV : _zz_8_string = "RISCV    ";
      IsaType_LOONGARCH : _zz_8_string = "LOONGARCH";
      default : _zz_8_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_10)
      ArchRegType_GPR : _zz_10_string = "GPR  ";
      ArchRegType_FPR : _zz_10_string = "FPR  ";
      ArchRegType_CSR : _zz_10_string = "CSR  ";
      ArchRegType_LA_CF : _zz_10_string = "LA_CF";
      default : _zz_10_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_13)
      ArchRegType_GPR : _zz_13_string = "GPR  ";
      ArchRegType_FPR : _zz_13_string = "FPR  ";
      ArchRegType_CSR : _zz_13_string = "CSR  ";
      ArchRegType_LA_CF : _zz_13_string = "LA_CF";
      default : _zz_13_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_16)
      ArchRegType_GPR : _zz_16_string = "GPR  ";
      ArchRegType_FPR : _zz_16_string = "FPR  ";
      ArchRegType_CSR : _zz_16_string = "CSR  ";
      ArchRegType_LA_CF : _zz_16_string = "LA_CF";
      default : _zz_16_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_20)
      ImmUsageType_NONE : _zz_20_string = "NONE         ";
      ImmUsageType_SRC_ALU : _zz_20_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : _zz_20_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : _zz_20_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : _zz_20_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : _zz_20_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : _zz_20_string = "JUMP_OFFSET  ";
      default : _zz_20_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_25)
      LogicOp_NONE : _zz_25_string = "NONE ";
      LogicOp_AND_1 : _zz_25_string = "AND_1";
      LogicOp_OR_1 : _zz_25_string = "OR_1 ";
      LogicOp_XOR_1 : _zz_25_string = "XOR_1";
      default : _zz_25_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_35)
      MemAccessSize_B : _zz_35_string = "B";
      MemAccessSize_H : _zz_35_string = "H";
      MemAccessSize_W : _zz_35_string = "W";
      MemAccessSize_D : _zz_35_string = "D";
      default : _zz_35_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_46)
      BranchCondition_NUL : _zz_46_string = "NUL        ";
      BranchCondition_EQ : _zz_46_string = "EQ         ";
      BranchCondition_NE : _zz_46_string = "NE         ";
      BranchCondition_LT : _zz_46_string = "LT         ";
      BranchCondition_GE : _zz_46_string = "GE         ";
      BranchCondition_LTU : _zz_46_string = "LTU        ";
      BranchCondition_GEU : _zz_46_string = "GEU        ";
      BranchCondition_EQZ : _zz_46_string = "EQZ        ";
      BranchCondition_NEZ : _zz_46_string = "NEZ        ";
      BranchCondition_LTZ : _zz_46_string = "LTZ        ";
      BranchCondition_GEZ : _zz_46_string = "GEZ        ";
      BranchCondition_GTZ : _zz_46_string = "GTZ        ";
      BranchCondition_LEZ : _zz_46_string = "LEZ        ";
      BranchCondition_F_EQ : _zz_46_string = "F_EQ       ";
      BranchCondition_F_NE : _zz_46_string = "F_NE       ";
      BranchCondition_F_LT : _zz_46_string = "F_LT       ";
      BranchCondition_F_LE : _zz_46_string = "F_LE       ";
      BranchCondition_F_UN : _zz_46_string = "F_UN       ";
      BranchCondition_LA_CF_TRUE : _zz_46_string = "LA_CF_TRUE ";
      BranchCondition_LA_CF_FALSE : _zz_46_string = "LA_CF_FALSE";
      default : _zz_46_string = "???????????";
    endcase
  end
  always @(*) begin
    case(_zz_50)
      ArchRegType_GPR : _zz_50_string = "GPR  ";
      ArchRegType_FPR : _zz_50_string = "FPR  ";
      ArchRegType_CSR : _zz_50_string = "CSR  ";
      ArchRegType_LA_CF : _zz_50_string = "LA_CF";
      default : _zz_50_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_54)
      MemAccessSize_B : _zz_54_string = "B";
      MemAccessSize_H : _zz_54_string = "H";
      MemAccessSize_W : _zz_54_string = "W";
      MemAccessSize_D : _zz_54_string = "D";
      default : _zz_54_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_55)
      MemAccessSize_B : _zz_55_string = "B";
      MemAccessSize_H : _zz_55_string = "H";
      MemAccessSize_W : _zz_55_string = "W";
      MemAccessSize_D : _zz_55_string = "D";
      default : _zz_55_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_56)
      MemAccessSize_B : _zz_56_string = "B";
      MemAccessSize_H : _zz_56_string = "H";
      MemAccessSize_W : _zz_56_string = "W";
      MemAccessSize_D : _zz_56_string = "D";
      default : _zz_56_string = "?";
    endcase
  end
  always @(*) begin
    case(_zz_71)
      DecodeExCode_INVALID : _zz_71_string = "INVALID     ";
      DecodeExCode_FETCH_ERROR : _zz_71_string = "FETCH_ERROR ";
      DecodeExCode_DECODE_ERROR : _zz_71_string = "DECODE_ERROR";
      DecodeExCode_OK : _zz_71_string = "OK          ";
      default : _zz_71_string = "????????????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    if(slotWillAllocate_0) begin
      _zz_1 = 1'b1;
    end
  end

  assign _zz_io_allocate_0_ready = (_zz__zz_io_allocate_0_ready < 4'b1000);
  assign io_allocate_0_ready = _zz_io_allocate_0_ready;
  assign io_canAllocate_0 = _zz_io_allocate_0_ready;
  assign slotWillAllocate_0 = (io_allocate_0_valid && io_allocate_0_ready);
  assign io_allocate_0_robPtr = (tailPtr_reg + 4'b0000);
  assign numActuallyAllocatedThisCycle = _zz_numActuallyAllocatedThisCycle;
  assign _zz_canCommitFlags_0 = (headPtr_reg + 4'b0000);
  assign _zz_io_commit_0_entry_status_busy = _zz_canCommitFlags_0[2:0];
  assign _zz_io_commit_0_entry_status_done = _zz__zz_io_commit_0_entry_status_done;
  assign _zz_io_commit_0_entry_status_genBit = _zz__zz_io_commit_0_entry_status_genBit;
  assign canCommitFlags_0 = ((((! ((io_flush_valid || flushInProgressReg) || flushWasActiveLastCycle)) && (4'b0000 < count_reg)) && _zz_io_commit_0_entry_status_done) && (_zz_canCommitFlags_0[3] == _zz_io_commit_0_entry_status_genBit));
  assign io_commit_0_valid = (4'b0000 < count_reg);
  assign io_commit_0_canCommit = canCommitFlags_0;
  assign _zz_io_commit_0_entry_payload_pc = payloads_spinal_port0;
  assign _zz_io_commit_0_entry_payload_uop_robPtr = _zz_io_commit_0_entry_payload_pc[337 : 0];
  assign _zz_io_commit_0_entry_payload_uop_decoded_pc = _zz_io_commit_0_entry_payload_uop_robPtr[276 : 0];
  assign _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1 = _zz_io_commit_0_entry_payload_uop_decoded_pc[37 : 33];
  assign _zz_io_commit_0_entry_payload_uop_decoded_uopCode = _zz_io_commit_0_entry_payload_uop_decoded_uopCode_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1 = _zz_io_commit_0_entry_payload_uop_decoded_pc[41 : 38];
  assign _zz_io_commit_0_entry_payload_uop_decoded_exeUnit = _zz_io_commit_0_entry_payload_uop_decoded_exeUnit_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_isa_1 = _zz_io_commit_0_entry_payload_uop_decoded_pc[43 : 42];
  assign _zz_io_commit_0_entry_payload_uop_decoded_isa = _zz_io_commit_0_entry_payload_uop_decoded_isa_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_archDest_idx = _zz_io_commit_0_entry_payload_uop_decoded_pc[50 : 44];
  assign _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1 = _zz_io_commit_0_entry_payload_uop_decoded_archDest_idx[6 : 5];
  assign _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype = _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_idx = _zz_io_commit_0_entry_payload_uop_decoded_pc[58 : 52];
  assign _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1 = _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_idx[6 : 5];
  assign _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype = _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_idx = _zz_io_commit_0_entry_payload_uop_decoded_pc[66 : 60];
  assign _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1 = _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_idx[6 : 5];
  assign _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype = _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1 = _zz_io_commit_0_entry_payload_uop_decoded_pc[103 : 101];
  assign _zz_io_commit_0_entry_payload_uop_decoded_immUsage = _zz_io_commit_0_entry_payload_uop_decoded_immUsage_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid = _zz_io_commit_0_entry_payload_uop_decoded_pc[109 : 104];
  assign _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1 = _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid[5 : 4];
  assign _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp = _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid = _zz_io_commit_0_entry_payload_uop_decoded_pc[114 : 110];
  assign _zz_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid = _zz_io_commit_0_entry_payload_uop_decoded_pc[118 : 115];
  assign _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad = _zz_io_commit_0_entry_payload_uop_decoded_pc[145 : 119];
  assign _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1 = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[1 : 0];
  assign _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump = _zz_io_commit_0_entry_payload_uop_decoded_pc[163 : 146];
  assign _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1 = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump[4 : 0];
  assign _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump[13 : 7];
  assign _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1 = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx[6 : 5];
  assign _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType = _zz_io_commit_0_entry_payload_uop_decoded_pc[184 : 164];
  assign _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1 = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[5 : 4];
  assign _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1 = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[7 : 6];
  assign _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1 = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[9 : 8];
  assign _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr = _zz_io_commit_0_entry_payload_uop_decoded_pc[202 : 185];
  assign _zz_io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode = _zz_io_commit_0_entry_payload_uop_decoded_pc[228 : 203];
  assign _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1 = _zz_io_commit_0_entry_payload_uop_decoded_pc[230 : 229];
  assign _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode = _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode_1;
  assign _zz_io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken = _zz_io_commit_0_entry_payload_uop_decoded_pc[276 : 243];
  assign _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx = _zz_io_commit_0_entry_payload_uop_robPtr[306 : 277];
  assign io_commit_0_entry_payload_uop_decoded_pc = _zz_io_commit_0_entry_payload_uop_decoded_pc[31 : 0];
  assign io_commit_0_entry_payload_uop_decoded_isValid = _zz_io_commit_0_entry_payload_uop_decoded_pc[32];
  assign io_commit_0_entry_payload_uop_decoded_uopCode = _zz_io_commit_0_entry_payload_uop_decoded_uopCode;
  assign io_commit_0_entry_payload_uop_decoded_exeUnit = _zz_io_commit_0_entry_payload_uop_decoded_exeUnit;
  assign io_commit_0_entry_payload_uop_decoded_isa = _zz_io_commit_0_entry_payload_uop_decoded_isa;
  assign io_commit_0_entry_payload_uop_decoded_archDest_idx = _zz_io_commit_0_entry_payload_uop_decoded_archDest_idx[4 : 0];
  assign io_commit_0_entry_payload_uop_decoded_archDest_rtype = _zz_io_commit_0_entry_payload_uop_decoded_archDest_rtype;
  assign io_commit_0_entry_payload_uop_decoded_writeArchDestEn = _zz_io_commit_0_entry_payload_uop_decoded_pc[51];
  assign io_commit_0_entry_payload_uop_decoded_archSrc1_idx = _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_idx[4 : 0];
  assign io_commit_0_entry_payload_uop_decoded_archSrc1_rtype = _zz_io_commit_0_entry_payload_uop_decoded_archSrc1_rtype;
  assign io_commit_0_entry_payload_uop_decoded_useArchSrc1 = _zz_io_commit_0_entry_payload_uop_decoded_pc[59];
  assign io_commit_0_entry_payload_uop_decoded_archSrc2_idx = _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_idx[4 : 0];
  assign io_commit_0_entry_payload_uop_decoded_archSrc2_rtype = _zz_io_commit_0_entry_payload_uop_decoded_archSrc2_rtype;
  assign io_commit_0_entry_payload_uop_decoded_useArchSrc2 = _zz_io_commit_0_entry_payload_uop_decoded_pc[67];
  assign io_commit_0_entry_payload_uop_decoded_usePcForAddr = _zz_io_commit_0_entry_payload_uop_decoded_pc[68];
  assign io_commit_0_entry_payload_uop_decoded_imm = _zz_io_commit_0_entry_payload_uop_decoded_pc[100 : 69];
  assign io_commit_0_entry_payload_uop_decoded_immUsage = _zz_io_commit_0_entry_payload_uop_decoded_immUsage;
  assign io_commit_0_entry_payload_uop_decoded_aluCtrl_valid = _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid[0];
  assign io_commit_0_entry_payload_uop_decoded_aluCtrl_isSub = _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid[1];
  assign io_commit_0_entry_payload_uop_decoded_aluCtrl_isAdd = _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid[2];
  assign io_commit_0_entry_payload_uop_decoded_aluCtrl_isSigned = _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_valid[3];
  assign io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp = _zz_io_commit_0_entry_payload_uop_decoded_aluCtrl_logicOp;
  assign io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid = _zz_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid[0];
  assign io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRight = _zz_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid[1];
  assign io_commit_0_entry_payload_uop_decoded_shiftCtrl_isArithmetic = _zz_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid[2];
  assign io_commit_0_entry_payload_uop_decoded_shiftCtrl_isRotate = _zz_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid[3];
  assign io_commit_0_entry_payload_uop_decoded_shiftCtrl_isDoubleWord = _zz_io_commit_0_entry_payload_uop_decoded_shiftCtrl_valid[4];
  assign io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid = _zz_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid[0];
  assign io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isDiv = _zz_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid[1];
  assign io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isSigned = _zz_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid[2];
  assign io_commit_0_entry_payload_uop_decoded_mulDivCtrl_isWordOp = _zz_io_commit_0_entry_payload_uop_decoded_mulDivCtrl_valid[3];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_size = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_size;
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[2];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_isStore = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[3];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_isLoadLinked = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[4];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_isStoreCond = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[5];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_atomicOp = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[10 : 6];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_isFence = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[11];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_fenceMode = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[19 : 12];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_isCacheOp = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[20];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_cacheOpType = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[25 : 21];
  assign io_commit_0_entry_payload_uop_decoded_memCtrl_isPrefetch = _zz_io_commit_0_entry_payload_uop_decoded_memCtrl_isSignedLoad[26];
  assign io_commit_0_entry_payload_uop_decoded_branchCtrl_condition = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_condition;
  assign io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump[5];
  assign io_commit_0_entry_payload_uop_decoded_branchCtrl_isLink = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump[6];
  assign io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_idx[4 : 0];
  assign io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_linkReg_rtype;
  assign io_commit_0_entry_payload_uop_decoded_branchCtrl_isIndirect = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump[14];
  assign io_commit_0_entry_payload_uop_decoded_branchCtrl_laCfIdx = _zz_io_commit_0_entry_payload_uop_decoded_branchCtrl_isJump[17 : 15];
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[3 : 0];
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1 = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc1;
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2 = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeSrc2;
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_fpSizeDest;
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_roundingMode = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[12 : 10];
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_isIntegerDest = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[13];
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_isSignedCvt = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[14];
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_fmaNegSrc1 = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[15];
  assign io_commit_0_entry_payload_uop_decoded_fpuCtrl_fcmpCond = _zz_io_commit_0_entry_payload_uop_decoded_fpuCtrl_opType[20 : 16];
  assign io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr = _zz_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr[13 : 0];
  assign io_commit_0_entry_payload_uop_decoded_csrCtrl_isWrite = _zz_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr[14];
  assign io_commit_0_entry_payload_uop_decoded_csrCtrl_isRead = _zz_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr[15];
  assign io_commit_0_entry_payload_uop_decoded_csrCtrl_isExchange = _zz_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr[16];
  assign io_commit_0_entry_payload_uop_decoded_csrCtrl_useUimmAsSrc = _zz_io_commit_0_entry_payload_uop_decoded_csrCtrl_csrAddr[17];
  assign io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode = _zz_io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode[19 : 0];
  assign io_commit_0_entry_payload_uop_decoded_sysCtrl_isExceptionReturn = _zz_io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode[20];
  assign io_commit_0_entry_payload_uop_decoded_sysCtrl_isTlbOp = _zz_io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode[21];
  assign io_commit_0_entry_payload_uop_decoded_sysCtrl_tlbOpType = _zz_io_commit_0_entry_payload_uop_decoded_sysCtrl_sysCode[25 : 22];
  assign io_commit_0_entry_payload_uop_decoded_decodeExceptionCode = _zz_io_commit_0_entry_payload_uop_decoded_decodeExceptionCode;
  assign io_commit_0_entry_payload_uop_decoded_hasDecodeException = _zz_io_commit_0_entry_payload_uop_decoded_pc[231];
  assign io_commit_0_entry_payload_uop_decoded_isMicrocode = _zz_io_commit_0_entry_payload_uop_decoded_pc[232];
  assign io_commit_0_entry_payload_uop_decoded_microcodeEntry = _zz_io_commit_0_entry_payload_uop_decoded_pc[240 : 233];
  assign io_commit_0_entry_payload_uop_decoded_isSerializing = _zz_io_commit_0_entry_payload_uop_decoded_pc[241];
  assign io_commit_0_entry_payload_uop_decoded_isBranchOrJump = _zz_io_commit_0_entry_payload_uop_decoded_pc[242];
  assign io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken = _zz_io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken[0];
  assign io_commit_0_entry_payload_uop_decoded_branchPrediction_target = _zz_io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken[32 : 1];
  assign io_commit_0_entry_payload_uop_decoded_branchPrediction_wasPredicted = _zz_io_commit_0_entry_payload_uop_decoded_branchPrediction_isTaken[33];
  assign io_commit_0_entry_payload_uop_rename_physSrc1_idx = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx_1[5 : 0];
  assign io_commit_0_entry_payload_uop_rename_physSrc1IsFpr = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[6];
  assign io_commit_0_entry_payload_uop_rename_physSrc2_idx = _zz_io_commit_0_entry_payload_uop_rename_physSrc2_idx[5 : 0];
  assign io_commit_0_entry_payload_uop_rename_physSrc2IsFpr = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[13];
  assign io_commit_0_entry_payload_uop_rename_physDest_idx = _zz_io_commit_0_entry_payload_uop_rename_physDest_idx[5 : 0];
  assign io_commit_0_entry_payload_uop_rename_physDestIsFpr = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[20];
  assign io_commit_0_entry_payload_uop_rename_oldPhysDest_idx = _zz_io_commit_0_entry_payload_uop_rename_oldPhysDest_idx[5 : 0];
  assign io_commit_0_entry_payload_uop_rename_oldPhysDestIsFpr = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[27];
  assign io_commit_0_entry_payload_uop_rename_allocatesPhysDest = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[28];
  assign io_commit_0_entry_payload_uop_rename_writesToPhysReg = _zz_io_commit_0_entry_payload_uop_rename_physSrc1_idx[29];
  assign io_commit_0_entry_payload_uop_robPtr = _zz_io_commit_0_entry_payload_uop_robPtr[310 : 307];
  assign io_commit_0_entry_payload_uop_uniqueId = _zz_io_commit_0_entry_payload_uop_robPtr[326 : 311];
  assign io_commit_0_entry_payload_uop_dispatched = _zz_io_commit_0_entry_payload_uop_robPtr[327];
  assign io_commit_0_entry_payload_uop_executed = _zz_io_commit_0_entry_payload_uop_robPtr[328];
  assign io_commit_0_entry_payload_uop_hasException = _zz_io_commit_0_entry_payload_uop_robPtr[329];
  assign io_commit_0_entry_payload_uop_exceptionCode = _zz_io_commit_0_entry_payload_uop_robPtr[337 : 330];
  assign io_commit_0_entry_payload_pc = _zz_io_commit_0_entry_payload_pc[369 : 338];
  assign io_commit_0_entry_status_busy = _zz_io_commit_0_entry_status_busy_1;
  assign io_commit_0_entry_status_done = _zz_io_commit_0_entry_status_done;
  assign io_commit_0_entry_status_isMispredictedBranch = _zz_io_commit_0_entry_status_isMispredictedBranch;
  assign io_commit_0_entry_status_isTaken = _zz_io_commit_0_entry_status_isTaken;
  assign io_commit_0_entry_status_result = _zz_io_commit_0_entry_status_result;
  assign io_commit_0_entry_status_hasException = _zz_io_commit_0_entry_status_hasException;
  assign io_commit_0_entry_status_exceptionCode = _zz_io_commit_0_entry_status_exceptionCode;
  assign io_commit_0_entry_status_genBit = _zz_io_commit_0_entry_status_genBit;
  assign actualCommittedMask_0 = ((1'b1 && canCommitFlags_0) && io_commitAck_0);
  assign numToCommit = _zz_numToCommit;
  assign when_ReorderBuffer_l285 = (1'b0 < numToCommit);
  always @(*) begin
    nextHead = (headPtr_reg + _zz_nextHead);
    if(io_flush_valid) begin
      case(io_flush_payload_reason)
        FlushReason_FULL_FLUSH : begin
          nextHead = 4'b0000;
        end
        FlushReason_ROLLBACK_TO_ROB_IDX : begin
          nextHead = headPtr_reg;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    nextTail = (tailPtr_reg + _zz_nextTail);
    if(io_flush_valid) begin
      case(io_flush_payload_reason)
        FlushReason_FULL_FLUSH : begin
          nextTail = 4'b0000;
        end
        FlushReason_ROLLBACK_TO_ROB_IDX : begin
          nextTail = io_flush_payload_targetRobPtr;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    nextCount = (_zz_nextCount_1 - _zz_nextCount_3);
    if(io_flush_valid) begin
      case(io_flush_payload_reason)
        FlushReason_FULL_FLUSH : begin
          nextCount = 4'b0000;
        end
        FlushReason_ROLLBACK_TO_ROB_IDX : begin
          nextCount = _zz_nextCount[3:0];
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_flushed = 1'b0;
    if(io_flush_valid) begin
      io_flushed = 1'b1;
    end
  end

  assign _zz_when_ReorderBuffer_l321 = {1'd0, headPtr_reg};
  assign _zz_when_ReorderBuffer_l321_1 = {1'd0, io_flush_payload_targetRobPtr};
  assign when_ReorderBuffer_l321 = (_zz_when_ReorderBuffer_l321 <= _zz_when_ReorderBuffer_l321_1);
  always @(*) begin
    if(when_ReorderBuffer_l321) begin
      _zz_nextCount = (_zz_when_ReorderBuffer_l321_1 - _zz_when_ReorderBuffer_l321);
    end else begin
      _zz_nextCount = (_zz__zz_nextCount + _zz__zz_nextCount_1);
    end
  end

  assign _zz_statuses_0_genBit = (tailPtr_reg + 4'b0000);
  assign _zz_3 = _zz_statuses_0_genBit[2:0];
  assign _zz_statuses_0_genBit_1 = _zz_statuses_0_genBit[3];
  assign _zz_4 = io_allocate_0_uopIn_decoded_pc;
  assign _zz_5 = io_allocate_0_uopIn_decoded_isValid;
  assign _zz_6 = io_allocate_0_uopIn_decoded_uopCode;
  assign _zz_7 = io_allocate_0_uopIn_decoded_exeUnit;
  assign _zz_8 = io_allocate_0_uopIn_decoded_isa;
  assign _zz_9 = io_allocate_0_uopIn_decoded_archDest_idx;
  assign _zz_10 = io_allocate_0_uopIn_decoded_archDest_rtype;
  assign _zz_11 = io_allocate_0_uopIn_decoded_writeArchDestEn;
  assign _zz_12 = io_allocate_0_uopIn_decoded_archSrc1_idx;
  assign _zz_13 = io_allocate_0_uopIn_decoded_archSrc1_rtype;
  assign _zz_14 = io_allocate_0_uopIn_decoded_useArchSrc1;
  assign _zz_15 = io_allocate_0_uopIn_decoded_archSrc2_idx;
  assign _zz_16 = io_allocate_0_uopIn_decoded_archSrc2_rtype;
  assign _zz_17 = io_allocate_0_uopIn_decoded_useArchSrc2;
  assign _zz_18 = io_allocate_0_uopIn_decoded_usePcForAddr;
  assign _zz_19 = io_allocate_0_uopIn_decoded_imm;
  assign _zz_20 = io_allocate_0_uopIn_decoded_immUsage;
  assign _zz_21 = io_allocate_0_uopIn_decoded_aluCtrl_valid;
  assign _zz_22 = io_allocate_0_uopIn_decoded_aluCtrl_isSub;
  assign _zz_23 = io_allocate_0_uopIn_decoded_aluCtrl_isAdd;
  assign _zz_24 = io_allocate_0_uopIn_decoded_aluCtrl_isSigned;
  assign _zz_25 = io_allocate_0_uopIn_decoded_aluCtrl_logicOp;
  assign _zz_26 = io_allocate_0_uopIn_decoded_shiftCtrl_valid;
  assign _zz_27 = io_allocate_0_uopIn_decoded_shiftCtrl_isRight;
  assign _zz_28 = io_allocate_0_uopIn_decoded_shiftCtrl_isArithmetic;
  assign _zz_29 = io_allocate_0_uopIn_decoded_shiftCtrl_isRotate;
  assign _zz_30 = io_allocate_0_uopIn_decoded_shiftCtrl_isDoubleWord;
  assign _zz_31 = io_allocate_0_uopIn_decoded_mulDivCtrl_valid;
  assign _zz_32 = io_allocate_0_uopIn_decoded_mulDivCtrl_isDiv;
  assign _zz_33 = io_allocate_0_uopIn_decoded_mulDivCtrl_isSigned;
  assign _zz_34 = io_allocate_0_uopIn_decoded_mulDivCtrl_isWordOp;
  assign _zz_35 = io_allocate_0_uopIn_decoded_memCtrl_size;
  assign _zz_36 = io_allocate_0_uopIn_decoded_memCtrl_isSignedLoad;
  assign _zz_37 = io_allocate_0_uopIn_decoded_memCtrl_isStore;
  assign _zz_38 = io_allocate_0_uopIn_decoded_memCtrl_isLoadLinked;
  assign _zz_39 = io_allocate_0_uopIn_decoded_memCtrl_isStoreCond;
  assign _zz_40 = io_allocate_0_uopIn_decoded_memCtrl_atomicOp;
  assign _zz_41 = io_allocate_0_uopIn_decoded_memCtrl_isFence;
  assign _zz_42 = io_allocate_0_uopIn_decoded_memCtrl_fenceMode;
  assign _zz_43 = io_allocate_0_uopIn_decoded_memCtrl_isCacheOp;
  assign _zz_44 = io_allocate_0_uopIn_decoded_memCtrl_cacheOpType;
  assign _zz_45 = io_allocate_0_uopIn_decoded_memCtrl_isPrefetch;
  assign _zz_46 = io_allocate_0_uopIn_decoded_branchCtrl_condition;
  assign _zz_47 = io_allocate_0_uopIn_decoded_branchCtrl_isJump;
  assign _zz_48 = io_allocate_0_uopIn_decoded_branchCtrl_isLink;
  assign _zz_49 = io_allocate_0_uopIn_decoded_branchCtrl_linkReg_idx;
  assign _zz_50 = io_allocate_0_uopIn_decoded_branchCtrl_linkReg_rtype;
  assign _zz_51 = io_allocate_0_uopIn_decoded_branchCtrl_isIndirect;
  assign _zz_52 = io_allocate_0_uopIn_decoded_branchCtrl_laCfIdx;
  assign _zz_53 = io_allocate_0_uopIn_decoded_fpuCtrl_opType;
  assign _zz_54 = io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc1;
  assign _zz_55 = io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeSrc2;
  assign _zz_56 = io_allocate_0_uopIn_decoded_fpuCtrl_fpSizeDest;
  assign _zz_57 = io_allocate_0_uopIn_decoded_fpuCtrl_roundingMode;
  assign _zz_58 = io_allocate_0_uopIn_decoded_fpuCtrl_isIntegerDest;
  assign _zz_59 = io_allocate_0_uopIn_decoded_fpuCtrl_isSignedCvt;
  assign _zz_60 = io_allocate_0_uopIn_decoded_fpuCtrl_fmaNegSrc1;
  assign _zz_61 = io_allocate_0_uopIn_decoded_fpuCtrl_fcmpCond;
  assign _zz_62 = io_allocate_0_uopIn_decoded_csrCtrl_csrAddr;
  assign _zz_63 = io_allocate_0_uopIn_decoded_csrCtrl_isWrite;
  assign _zz_64 = io_allocate_0_uopIn_decoded_csrCtrl_isRead;
  assign _zz_65 = io_allocate_0_uopIn_decoded_csrCtrl_isExchange;
  assign _zz_66 = io_allocate_0_uopIn_decoded_csrCtrl_useUimmAsSrc;
  assign _zz_67 = io_allocate_0_uopIn_decoded_sysCtrl_sysCode;
  assign _zz_68 = io_allocate_0_uopIn_decoded_sysCtrl_isExceptionReturn;
  assign _zz_69 = io_allocate_0_uopIn_decoded_sysCtrl_isTlbOp;
  assign _zz_70 = io_allocate_0_uopIn_decoded_sysCtrl_tlbOpType;
  assign _zz_71 = io_allocate_0_uopIn_decoded_decodeExceptionCode;
  assign _zz_72 = io_allocate_0_uopIn_decoded_hasDecodeException;
  assign _zz_73 = io_allocate_0_uopIn_decoded_isMicrocode;
  assign _zz_74 = io_allocate_0_uopIn_decoded_microcodeEntry;
  assign _zz_75 = io_allocate_0_uopIn_decoded_isSerializing;
  assign _zz_76 = io_allocate_0_uopIn_decoded_isBranchOrJump;
  assign _zz_77 = io_allocate_0_uopIn_decoded_branchPrediction_isTaken;
  assign _zz_78 = io_allocate_0_uopIn_decoded_branchPrediction_target;
  assign _zz_79 = io_allocate_0_uopIn_decoded_branchPrediction_wasPredicted;
  assign _zz_80 = io_allocate_0_uopIn_rename_physSrc1_idx;
  assign _zz_81 = io_allocate_0_uopIn_rename_physSrc1IsFpr;
  assign _zz_82 = io_allocate_0_uopIn_rename_physSrc2_idx;
  assign _zz_83 = io_allocate_0_uopIn_rename_physSrc2IsFpr;
  assign _zz_84 = io_allocate_0_uopIn_rename_physDest_idx;
  assign _zz_85 = io_allocate_0_uopIn_rename_physDestIsFpr;
  assign _zz_86 = io_allocate_0_uopIn_rename_oldPhysDest_idx;
  assign _zz_87 = io_allocate_0_uopIn_rename_oldPhysDestIsFpr;
  assign _zz_88 = io_allocate_0_uopIn_rename_allocatesPhysDest;
  assign _zz_89 = io_allocate_0_uopIn_rename_writesToPhysReg;
  always @(*) begin
    _zz_90 = io_allocate_0_uopIn_robPtr;
    _zz_90 = _zz_statuses_0_genBit;
  end

  assign _zz_91 = io_allocate_0_uopIn_uniqueId;
  assign _zz_92 = io_allocate_0_uopIn_dispatched;
  assign _zz_93 = io_allocate_0_uopIn_executed;
  assign _zz_94 = io_allocate_0_uopIn_hasException;
  assign _zz_95 = io_allocate_0_uopIn_exceptionCode;
  assign _zz_96 = io_allocate_0_pcIn;
  assign _zz_97 = ({7'd0,1'b1} <<< _zz_3);
  assign _zz_98 = _zz_97[0];
  assign _zz_99 = _zz_97[1];
  assign _zz_100 = _zz_97[2];
  assign _zz_101 = _zz_97[3];
  assign _zz_102 = _zz_97[4];
  assign _zz_103 = _zz_97[5];
  assign _zz_104 = _zz_97[6];
  assign _zz_105 = _zz_97[7];
  assign _zz_when_ReorderBuffer_l375 = io_writeback_0_robPtr[2:0];
  assign _zz_107 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l375);
  assign _zz_108 = _zz_107[0];
  assign _zz_109 = _zz_107[1];
  assign _zz_110 = _zz_107[2];
  assign _zz_111 = _zz_107[3];
  assign _zz_112 = _zz_107[4];
  assign _zz_113 = _zz_107[5];
  assign _zz_114 = _zz_107[6];
  assign _zz_115 = _zz_107[7];
  assign when_ReorderBuffer_l375 = (((! io_flush_valid) && io_writeback_0_fire) && (io_writeback_0_robPtr[3] == _zz_when_ReorderBuffer_l375_5));
  assign _zz_statuses_0_exceptionCode = (io_writeback_0_exceptionOccurred ? io_writeback_0_exceptionCodeIn : _zz__zz_statuses_0_exceptionCode);
  assign _zz_when_ReorderBuffer_l375_1 = io_writeback_1_robPtr[2:0];
  assign _zz_116 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l375_1);
  assign _zz_117 = _zz_116[0];
  assign _zz_118 = _zz_116[1];
  assign _zz_119 = _zz_116[2];
  assign _zz_120 = _zz_116[3];
  assign _zz_121 = _zz_116[4];
  assign _zz_122 = _zz_116[5];
  assign _zz_123 = _zz_116[6];
  assign _zz_124 = _zz_116[7];
  assign when_ReorderBuffer_l375_1 = (((! io_flush_valid) && io_writeback_1_fire) && (io_writeback_1_robPtr[3] == _zz_when_ReorderBuffer_l375_1_1));
  assign _zz_statuses_0_exceptionCode_1 = (io_writeback_1_exceptionOccurred ? io_writeback_1_exceptionCodeIn : _zz__zz_statuses_0_exceptionCode_1);
  assign _zz_when_ReorderBuffer_l375_2 = io_writeback_2_robPtr[2:0];
  assign _zz_125 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l375_2);
  assign _zz_126 = _zz_125[0];
  assign _zz_127 = _zz_125[1];
  assign _zz_128 = _zz_125[2];
  assign _zz_129 = _zz_125[3];
  assign _zz_130 = _zz_125[4];
  assign _zz_131 = _zz_125[5];
  assign _zz_132 = _zz_125[6];
  assign _zz_133 = _zz_125[7];
  assign when_ReorderBuffer_l375_2 = (((! io_flush_valid) && io_writeback_2_fire) && (io_writeback_2_robPtr[3] == _zz_when_ReorderBuffer_l375_2_1));
  assign _zz_statuses_0_exceptionCode_2 = (io_writeback_2_exceptionOccurred ? io_writeback_2_exceptionCodeIn : _zz__zz_statuses_0_exceptionCode_2);
  assign _zz_when_ReorderBuffer_l375_3 = io_writeback_3_robPtr[2:0];
  assign _zz_134 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l375_3);
  assign _zz_135 = _zz_134[0];
  assign _zz_136 = _zz_134[1];
  assign _zz_137 = _zz_134[2];
  assign _zz_138 = _zz_134[3];
  assign _zz_139 = _zz_134[4];
  assign _zz_140 = _zz_134[5];
  assign _zz_141 = _zz_134[6];
  assign _zz_142 = _zz_134[7];
  assign when_ReorderBuffer_l375_3 = (((! io_flush_valid) && io_writeback_3_fire) && (io_writeback_3_robPtr[3] == _zz_when_ReorderBuffer_l375_3_1));
  assign _zz_statuses_0_exceptionCode_3 = (io_writeback_3_exceptionOccurred ? io_writeback_3_exceptionCodeIn : _zz__zz_statuses_0_exceptionCode_3);
  assign _zz_when_ReorderBuffer_l375_4 = io_writeback_4_robPtr[2:0];
  assign _zz_143 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l375_4);
  assign _zz_144 = _zz_143[0];
  assign _zz_145 = _zz_143[1];
  assign _zz_146 = _zz_143[2];
  assign _zz_147 = _zz_143[3];
  assign _zz_148 = _zz_143[4];
  assign _zz_149 = _zz_143[5];
  assign _zz_150 = _zz_143[6];
  assign _zz_151 = _zz_143[7];
  assign when_ReorderBuffer_l375_4 = (((! io_flush_valid) && io_writeback_4_fire) && (io_writeback_4_robPtr[3] == _zz_when_ReorderBuffer_l375_4_1));
  assign _zz_statuses_0_exceptionCode_4 = (io_writeback_4_exceptionOccurred ? io_writeback_4_exceptionCodeIn : _zz__zz_statuses_0_exceptionCode_4);
  assign _zz_when_ReorderBuffer_l418 = 3'b000;
  assign _zz_152 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l418);
  assign _zz_153 = _zz_152[0];
  assign _zz_154 = _zz_152[1];
  assign _zz_155 = _zz_152[2];
  assign _zz_156 = _zz_152[3];
  assign _zz_157 = _zz_152[4];
  assign _zz_158 = _zz_152[5];
  assign _zz_159 = _zz_152[6];
  assign _zz_160 = _zz_152[7];
  assign _zz_when_ReorderBuffer_l418_1 = {1'd0, io_flush_payload_targetRobPtr};
  assign _zz_when_ReorderBuffer_l418_2 = {1'd0, tailPtr_reg};
  assign _zz_when_ReorderBuffer_l418_3 = {1'd0, _zz__zz_when_ReorderBuffer_l418_3};
  assign when_ReorderBuffer_l412 = (_zz_when_ReorderBuffer_l418_1 <= _zz_when_ReorderBuffer_l418_2);
  always @(*) begin
    if(when_ReorderBuffer_l412) begin
      when_ReorderBuffer_l418 = ((_zz_when_ReorderBuffer_l418_1 <= _zz_when_ReorderBuffer_l418_3) && (_zz_when_ReorderBuffer_l418_3 < _zz_when_ReorderBuffer_l418_2));
    end else begin
      when_ReorderBuffer_l418 = ((_zz_when_ReorderBuffer_l418_1 <= _zz_when_ReorderBuffer_l418_3) || (_zz_when_ReorderBuffer_l418_3 < _zz_when_ReorderBuffer_l418_2));
    end
  end

  assign _zz_when_ReorderBuffer_l418_4 = 3'b001;
  assign _zz_161 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l418_4);
  assign _zz_162 = _zz_161[0];
  assign _zz_163 = _zz_161[1];
  assign _zz_164 = _zz_161[2];
  assign _zz_165 = _zz_161[3];
  assign _zz_166 = _zz_161[4];
  assign _zz_167 = _zz_161[5];
  assign _zz_168 = _zz_161[6];
  assign _zz_169 = _zz_161[7];
  assign _zz_when_ReorderBuffer_l418_5 = {1'd0, io_flush_payload_targetRobPtr};
  assign _zz_when_ReorderBuffer_l418_6 = {1'd0, tailPtr_reg};
  assign _zz_when_ReorderBuffer_l418_7 = {1'd0, _zz__zz_when_ReorderBuffer_l418_7};
  assign when_ReorderBuffer_l412_1 = (_zz_when_ReorderBuffer_l418_5 <= _zz_when_ReorderBuffer_l418_6);
  always @(*) begin
    if(when_ReorderBuffer_l412_1) begin
      when_ReorderBuffer_l418_1 = ((_zz_when_ReorderBuffer_l418_5 <= _zz_when_ReorderBuffer_l418_7) && (_zz_when_ReorderBuffer_l418_7 < _zz_when_ReorderBuffer_l418_6));
    end else begin
      when_ReorderBuffer_l418_1 = ((_zz_when_ReorderBuffer_l418_5 <= _zz_when_ReorderBuffer_l418_7) || (_zz_when_ReorderBuffer_l418_7 < _zz_when_ReorderBuffer_l418_6));
    end
  end

  assign _zz_when_ReorderBuffer_l418_8 = 3'b010;
  assign _zz_170 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l418_8);
  assign _zz_171 = _zz_170[0];
  assign _zz_172 = _zz_170[1];
  assign _zz_173 = _zz_170[2];
  assign _zz_174 = _zz_170[3];
  assign _zz_175 = _zz_170[4];
  assign _zz_176 = _zz_170[5];
  assign _zz_177 = _zz_170[6];
  assign _zz_178 = _zz_170[7];
  assign _zz_when_ReorderBuffer_l418_9 = {1'd0, io_flush_payload_targetRobPtr};
  assign _zz_when_ReorderBuffer_l418_10 = {1'd0, tailPtr_reg};
  assign _zz_when_ReorderBuffer_l418_11 = {1'd0, _zz__zz_when_ReorderBuffer_l418_11};
  assign when_ReorderBuffer_l412_2 = (_zz_when_ReorderBuffer_l418_9 <= _zz_when_ReorderBuffer_l418_10);
  always @(*) begin
    if(when_ReorderBuffer_l412_2) begin
      when_ReorderBuffer_l418_2 = ((_zz_when_ReorderBuffer_l418_9 <= _zz_when_ReorderBuffer_l418_11) && (_zz_when_ReorderBuffer_l418_11 < _zz_when_ReorderBuffer_l418_10));
    end else begin
      when_ReorderBuffer_l418_2 = ((_zz_when_ReorderBuffer_l418_9 <= _zz_when_ReorderBuffer_l418_11) || (_zz_when_ReorderBuffer_l418_11 < _zz_when_ReorderBuffer_l418_10));
    end
  end

  assign _zz_when_ReorderBuffer_l418_12 = 3'b011;
  assign _zz_179 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l418_12);
  assign _zz_180 = _zz_179[0];
  assign _zz_181 = _zz_179[1];
  assign _zz_182 = _zz_179[2];
  assign _zz_183 = _zz_179[3];
  assign _zz_184 = _zz_179[4];
  assign _zz_185 = _zz_179[5];
  assign _zz_186 = _zz_179[6];
  assign _zz_187 = _zz_179[7];
  assign _zz_when_ReorderBuffer_l418_13 = {1'd0, io_flush_payload_targetRobPtr};
  assign _zz_when_ReorderBuffer_l418_14 = {1'd0, tailPtr_reg};
  assign _zz_when_ReorderBuffer_l418_15 = {1'd0, _zz__zz_when_ReorderBuffer_l418_15};
  assign when_ReorderBuffer_l412_3 = (_zz_when_ReorderBuffer_l418_13 <= _zz_when_ReorderBuffer_l418_14);
  always @(*) begin
    if(when_ReorderBuffer_l412_3) begin
      when_ReorderBuffer_l418_3 = ((_zz_when_ReorderBuffer_l418_13 <= _zz_when_ReorderBuffer_l418_15) && (_zz_when_ReorderBuffer_l418_15 < _zz_when_ReorderBuffer_l418_14));
    end else begin
      when_ReorderBuffer_l418_3 = ((_zz_when_ReorderBuffer_l418_13 <= _zz_when_ReorderBuffer_l418_15) || (_zz_when_ReorderBuffer_l418_15 < _zz_when_ReorderBuffer_l418_14));
    end
  end

  assign _zz_when_ReorderBuffer_l418_16 = 3'b100;
  assign _zz_188 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l418_16);
  assign _zz_189 = _zz_188[0];
  assign _zz_190 = _zz_188[1];
  assign _zz_191 = _zz_188[2];
  assign _zz_192 = _zz_188[3];
  assign _zz_193 = _zz_188[4];
  assign _zz_194 = _zz_188[5];
  assign _zz_195 = _zz_188[6];
  assign _zz_196 = _zz_188[7];
  assign _zz_when_ReorderBuffer_l418_17 = {1'd0, io_flush_payload_targetRobPtr};
  assign _zz_when_ReorderBuffer_l418_18 = {1'd0, tailPtr_reg};
  assign _zz_when_ReorderBuffer_l418_19 = {1'd0, _zz__zz_when_ReorderBuffer_l418_19};
  assign when_ReorderBuffer_l412_4 = (_zz_when_ReorderBuffer_l418_17 <= _zz_when_ReorderBuffer_l418_18);
  always @(*) begin
    if(when_ReorderBuffer_l412_4) begin
      when_ReorderBuffer_l418_4 = ((_zz_when_ReorderBuffer_l418_17 <= _zz_when_ReorderBuffer_l418_19) && (_zz_when_ReorderBuffer_l418_19 < _zz_when_ReorderBuffer_l418_18));
    end else begin
      when_ReorderBuffer_l418_4 = ((_zz_when_ReorderBuffer_l418_17 <= _zz_when_ReorderBuffer_l418_19) || (_zz_when_ReorderBuffer_l418_19 < _zz_when_ReorderBuffer_l418_18));
    end
  end

  assign _zz_when_ReorderBuffer_l418_20 = 3'b101;
  assign _zz_197 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l418_20);
  assign _zz_198 = _zz_197[0];
  assign _zz_199 = _zz_197[1];
  assign _zz_200 = _zz_197[2];
  assign _zz_201 = _zz_197[3];
  assign _zz_202 = _zz_197[4];
  assign _zz_203 = _zz_197[5];
  assign _zz_204 = _zz_197[6];
  assign _zz_205 = _zz_197[7];
  assign _zz_when_ReorderBuffer_l418_21 = {1'd0, io_flush_payload_targetRobPtr};
  assign _zz_when_ReorderBuffer_l418_22 = {1'd0, tailPtr_reg};
  assign _zz_when_ReorderBuffer_l418_23 = {1'd0, _zz__zz_when_ReorderBuffer_l418_23};
  assign when_ReorderBuffer_l412_5 = (_zz_when_ReorderBuffer_l418_21 <= _zz_when_ReorderBuffer_l418_22);
  always @(*) begin
    if(when_ReorderBuffer_l412_5) begin
      when_ReorderBuffer_l418_5 = ((_zz_when_ReorderBuffer_l418_21 <= _zz_when_ReorderBuffer_l418_23) && (_zz_when_ReorderBuffer_l418_23 < _zz_when_ReorderBuffer_l418_22));
    end else begin
      when_ReorderBuffer_l418_5 = ((_zz_when_ReorderBuffer_l418_21 <= _zz_when_ReorderBuffer_l418_23) || (_zz_when_ReorderBuffer_l418_23 < _zz_when_ReorderBuffer_l418_22));
    end
  end

  assign _zz_when_ReorderBuffer_l418_24 = 3'b110;
  assign _zz_206 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l418_24);
  assign _zz_207 = _zz_206[0];
  assign _zz_208 = _zz_206[1];
  assign _zz_209 = _zz_206[2];
  assign _zz_210 = _zz_206[3];
  assign _zz_211 = _zz_206[4];
  assign _zz_212 = _zz_206[5];
  assign _zz_213 = _zz_206[6];
  assign _zz_214 = _zz_206[7];
  assign _zz_when_ReorderBuffer_l418_25 = {1'd0, io_flush_payload_targetRobPtr};
  assign _zz_when_ReorderBuffer_l418_26 = {1'd0, tailPtr_reg};
  assign _zz_when_ReorderBuffer_l418_27 = {1'd0, _zz__zz_when_ReorderBuffer_l418_27};
  assign when_ReorderBuffer_l412_6 = (_zz_when_ReorderBuffer_l418_25 <= _zz_when_ReorderBuffer_l418_26);
  always @(*) begin
    if(when_ReorderBuffer_l412_6) begin
      when_ReorderBuffer_l418_6 = ((_zz_when_ReorderBuffer_l418_25 <= _zz_when_ReorderBuffer_l418_27) && (_zz_when_ReorderBuffer_l418_27 < _zz_when_ReorderBuffer_l418_26));
    end else begin
      when_ReorderBuffer_l418_6 = ((_zz_when_ReorderBuffer_l418_25 <= _zz_when_ReorderBuffer_l418_27) || (_zz_when_ReorderBuffer_l418_27 < _zz_when_ReorderBuffer_l418_26));
    end
  end

  assign _zz_when_ReorderBuffer_l418_28 = 3'b111;
  assign _zz_215 = ({7'd0,1'b1} <<< _zz_when_ReorderBuffer_l418_28);
  assign _zz_216 = _zz_215[0];
  assign _zz_217 = _zz_215[1];
  assign _zz_218 = _zz_215[2];
  assign _zz_219 = _zz_215[3];
  assign _zz_220 = _zz_215[4];
  assign _zz_221 = _zz_215[5];
  assign _zz_222 = _zz_215[6];
  assign _zz_223 = _zz_215[7];
  assign _zz_when_ReorderBuffer_l418_29 = {1'd0, io_flush_payload_targetRobPtr};
  assign _zz_when_ReorderBuffer_l418_30 = {1'd0, tailPtr_reg};
  assign _zz_when_ReorderBuffer_l418_31 = {1'd0, _zz__zz_when_ReorderBuffer_l418_31};
  assign when_ReorderBuffer_l412_7 = (_zz_when_ReorderBuffer_l418_29 <= _zz_when_ReorderBuffer_l418_30);
  always @(*) begin
    if(when_ReorderBuffer_l412_7) begin
      when_ReorderBuffer_l418_7 = ((_zz_when_ReorderBuffer_l418_29 <= _zz_when_ReorderBuffer_l418_31) && (_zz_when_ReorderBuffer_l418_31 < _zz_when_ReorderBuffer_l418_30));
    end else begin
      when_ReorderBuffer_l418_7 = ((_zz_when_ReorderBuffer_l418_29 <= _zz_when_ReorderBuffer_l418_31) || (_zz_when_ReorderBuffer_l418_31 < _zz_when_ReorderBuffer_l418_30));
    end
  end

  assign io_empty = (count_reg == 4'b0000);
  assign io_headPtrOut = headPtr_reg;
  assign io_tailPtrOut = tailPtr_reg;
  assign io_countOut = count_reg;
  always @(posedge clk) begin
    if(reset) begin
      statuses_0_busy <= 1'b0;
      statuses_0_done <= 1'b0;
      statuses_0_hasException <= 1'b0;
      statuses_0_exceptionCode <= 8'h0;
      statuses_0_genBit <= 1'b0;
      statuses_1_busy <= 1'b0;
      statuses_1_done <= 1'b0;
      statuses_1_hasException <= 1'b0;
      statuses_1_exceptionCode <= 8'h0;
      statuses_1_genBit <= 1'b0;
      statuses_2_busy <= 1'b0;
      statuses_2_done <= 1'b0;
      statuses_2_hasException <= 1'b0;
      statuses_2_exceptionCode <= 8'h0;
      statuses_2_genBit <= 1'b0;
      statuses_3_busy <= 1'b0;
      statuses_3_done <= 1'b0;
      statuses_3_hasException <= 1'b0;
      statuses_3_exceptionCode <= 8'h0;
      statuses_3_genBit <= 1'b0;
      statuses_4_busy <= 1'b0;
      statuses_4_done <= 1'b0;
      statuses_4_hasException <= 1'b0;
      statuses_4_exceptionCode <= 8'h0;
      statuses_4_genBit <= 1'b0;
      statuses_5_busy <= 1'b0;
      statuses_5_done <= 1'b0;
      statuses_5_hasException <= 1'b0;
      statuses_5_exceptionCode <= 8'h0;
      statuses_5_genBit <= 1'b0;
      statuses_6_busy <= 1'b0;
      statuses_6_done <= 1'b0;
      statuses_6_hasException <= 1'b0;
      statuses_6_exceptionCode <= 8'h0;
      statuses_6_genBit <= 1'b0;
      statuses_7_busy <= 1'b0;
      statuses_7_done <= 1'b0;
      statuses_7_hasException <= 1'b0;
      statuses_7_exceptionCode <= 8'h0;
      statuses_7_genBit <= 1'b0;
      headPtr_reg <= 4'b0000;
      tailPtr_reg <= 4'b0000;
      count_reg <= 4'b0000;
      flushInProgressReg <= 1'b0;
      flushWasActiveLastCycle <= 1'b0;
    end else begin
      flushWasActiveLastCycle <= io_flush_valid;
      if(io_flush_valid) begin
        flushInProgressReg <= 1'b1;
      end else begin
        if(flushWasActiveLastCycle) begin
          flushInProgressReg <= 1'b0;
        end
      end
      if(when_ReorderBuffer_l285) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // ReorderBuffer.scala:L286
          `else
            if(!1'b0) begin
              $display("NOTE(ReorderBuffer.scala:286):  [ROB] COMMIT_SUMMARY: Committing %x entries, total entries=%x, capacity=8", numToCommit, count_reg); // ReorderBuffer.scala:L286
            end
          `endif
        `endif
      end
      headPtr_reg <= nextHead;
      tailPtr_reg <= nextTail;
      count_reg <= nextCount;
      if(slotWillAllocate_0) begin
        if(_zz_98) begin
          statuses_0_busy <= 1'b1;
        end
        if(_zz_99) begin
          statuses_1_busy <= 1'b1;
        end
        if(_zz_100) begin
          statuses_2_busy <= 1'b1;
        end
        if(_zz_101) begin
          statuses_3_busy <= 1'b1;
        end
        if(_zz_102) begin
          statuses_4_busy <= 1'b1;
        end
        if(_zz_103) begin
          statuses_5_busy <= 1'b1;
        end
        if(_zz_104) begin
          statuses_6_busy <= 1'b1;
        end
        if(_zz_105) begin
          statuses_7_busy <= 1'b1;
        end
        if(_zz_98) begin
          statuses_0_done <= 1'b0;
        end
        if(_zz_99) begin
          statuses_1_done <= 1'b0;
        end
        if(_zz_100) begin
          statuses_2_done <= 1'b0;
        end
        if(_zz_101) begin
          statuses_3_done <= 1'b0;
        end
        if(_zz_102) begin
          statuses_4_done <= 1'b0;
        end
        if(_zz_103) begin
          statuses_5_done <= 1'b0;
        end
        if(_zz_104) begin
          statuses_6_done <= 1'b0;
        end
        if(_zz_105) begin
          statuses_7_done <= 1'b0;
        end
        if(_zz_98) begin
          statuses_0_hasException <= 1'b0;
        end
        if(_zz_99) begin
          statuses_1_hasException <= 1'b0;
        end
        if(_zz_100) begin
          statuses_2_hasException <= 1'b0;
        end
        if(_zz_101) begin
          statuses_3_hasException <= 1'b0;
        end
        if(_zz_102) begin
          statuses_4_hasException <= 1'b0;
        end
        if(_zz_103) begin
          statuses_5_hasException <= 1'b0;
        end
        if(_zz_104) begin
          statuses_6_hasException <= 1'b0;
        end
        if(_zz_105) begin
          statuses_7_hasException <= 1'b0;
        end
        if(_zz_98) begin
          statuses_0_genBit <= _zz_statuses_0_genBit_1;
        end
        if(_zz_99) begin
          statuses_1_genBit <= _zz_statuses_0_genBit_1;
        end
        if(_zz_100) begin
          statuses_2_genBit <= _zz_statuses_0_genBit_1;
        end
        if(_zz_101) begin
          statuses_3_genBit <= _zz_statuses_0_genBit_1;
        end
        if(_zz_102) begin
          statuses_4_genBit <= _zz_statuses_0_genBit_1;
        end
        if(_zz_103) begin
          statuses_5_genBit <= _zz_statuses_0_genBit_1;
        end
        if(_zz_104) begin
          statuses_6_genBit <= _zz_statuses_0_genBit_1;
        end
        if(_zz_105) begin
          statuses_7_genBit <= _zz_statuses_0_genBit_1;
        end
      end
      if(when_ReorderBuffer_l375) begin
        if(_zz_108) begin
          statuses_0_busy <= 1'b0;
        end
        if(_zz_109) begin
          statuses_1_busy <= 1'b0;
        end
        if(_zz_110) begin
          statuses_2_busy <= 1'b0;
        end
        if(_zz_111) begin
          statuses_3_busy <= 1'b0;
        end
        if(_zz_112) begin
          statuses_4_busy <= 1'b0;
        end
        if(_zz_113) begin
          statuses_5_busy <= 1'b0;
        end
        if(_zz_114) begin
          statuses_6_busy <= 1'b0;
        end
        if(_zz_115) begin
          statuses_7_busy <= 1'b0;
        end
        if(_zz_108) begin
          statuses_0_done <= 1'b1;
        end
        if(_zz_109) begin
          statuses_1_done <= 1'b1;
        end
        if(_zz_110) begin
          statuses_2_done <= 1'b1;
        end
        if(_zz_111) begin
          statuses_3_done <= 1'b1;
        end
        if(_zz_112) begin
          statuses_4_done <= 1'b1;
        end
        if(_zz_113) begin
          statuses_5_done <= 1'b1;
        end
        if(_zz_114) begin
          statuses_6_done <= 1'b1;
        end
        if(_zz_115) begin
          statuses_7_done <= 1'b1;
        end
        if(_zz_108) begin
          statuses_0_hasException <= io_writeback_0_exceptionOccurred;
        end
        if(_zz_109) begin
          statuses_1_hasException <= io_writeback_0_exceptionOccurred;
        end
        if(_zz_110) begin
          statuses_2_hasException <= io_writeback_0_exceptionOccurred;
        end
        if(_zz_111) begin
          statuses_3_hasException <= io_writeback_0_exceptionOccurred;
        end
        if(_zz_112) begin
          statuses_4_hasException <= io_writeback_0_exceptionOccurred;
        end
        if(_zz_113) begin
          statuses_5_hasException <= io_writeback_0_exceptionOccurred;
        end
        if(_zz_114) begin
          statuses_6_hasException <= io_writeback_0_exceptionOccurred;
        end
        if(_zz_115) begin
          statuses_7_hasException <= io_writeback_0_exceptionOccurred;
        end
        if(_zz_108) begin
          statuses_0_exceptionCode <= _zz_statuses_0_exceptionCode;
        end
        if(_zz_109) begin
          statuses_1_exceptionCode <= _zz_statuses_0_exceptionCode;
        end
        if(_zz_110) begin
          statuses_2_exceptionCode <= _zz_statuses_0_exceptionCode;
        end
        if(_zz_111) begin
          statuses_3_exceptionCode <= _zz_statuses_0_exceptionCode;
        end
        if(_zz_112) begin
          statuses_4_exceptionCode <= _zz_statuses_0_exceptionCode;
        end
        if(_zz_113) begin
          statuses_5_exceptionCode <= _zz_statuses_0_exceptionCode;
        end
        if(_zz_114) begin
          statuses_6_exceptionCode <= _zz_statuses_0_exceptionCode;
        end
        if(_zz_115) begin
          statuses_7_exceptionCode <= _zz_statuses_0_exceptionCode;
        end
      end
      if(when_ReorderBuffer_l375_1) begin
        if(_zz_117) begin
          statuses_0_busy <= 1'b0;
        end
        if(_zz_118) begin
          statuses_1_busy <= 1'b0;
        end
        if(_zz_119) begin
          statuses_2_busy <= 1'b0;
        end
        if(_zz_120) begin
          statuses_3_busy <= 1'b0;
        end
        if(_zz_121) begin
          statuses_4_busy <= 1'b0;
        end
        if(_zz_122) begin
          statuses_5_busy <= 1'b0;
        end
        if(_zz_123) begin
          statuses_6_busy <= 1'b0;
        end
        if(_zz_124) begin
          statuses_7_busy <= 1'b0;
        end
        if(_zz_117) begin
          statuses_0_done <= 1'b1;
        end
        if(_zz_118) begin
          statuses_1_done <= 1'b1;
        end
        if(_zz_119) begin
          statuses_2_done <= 1'b1;
        end
        if(_zz_120) begin
          statuses_3_done <= 1'b1;
        end
        if(_zz_121) begin
          statuses_4_done <= 1'b1;
        end
        if(_zz_122) begin
          statuses_5_done <= 1'b1;
        end
        if(_zz_123) begin
          statuses_6_done <= 1'b1;
        end
        if(_zz_124) begin
          statuses_7_done <= 1'b1;
        end
        if(_zz_117) begin
          statuses_0_hasException <= io_writeback_1_exceptionOccurred;
        end
        if(_zz_118) begin
          statuses_1_hasException <= io_writeback_1_exceptionOccurred;
        end
        if(_zz_119) begin
          statuses_2_hasException <= io_writeback_1_exceptionOccurred;
        end
        if(_zz_120) begin
          statuses_3_hasException <= io_writeback_1_exceptionOccurred;
        end
        if(_zz_121) begin
          statuses_4_hasException <= io_writeback_1_exceptionOccurred;
        end
        if(_zz_122) begin
          statuses_5_hasException <= io_writeback_1_exceptionOccurred;
        end
        if(_zz_123) begin
          statuses_6_hasException <= io_writeback_1_exceptionOccurred;
        end
        if(_zz_124) begin
          statuses_7_hasException <= io_writeback_1_exceptionOccurred;
        end
        if(_zz_117) begin
          statuses_0_exceptionCode <= _zz_statuses_0_exceptionCode_1;
        end
        if(_zz_118) begin
          statuses_1_exceptionCode <= _zz_statuses_0_exceptionCode_1;
        end
        if(_zz_119) begin
          statuses_2_exceptionCode <= _zz_statuses_0_exceptionCode_1;
        end
        if(_zz_120) begin
          statuses_3_exceptionCode <= _zz_statuses_0_exceptionCode_1;
        end
        if(_zz_121) begin
          statuses_4_exceptionCode <= _zz_statuses_0_exceptionCode_1;
        end
        if(_zz_122) begin
          statuses_5_exceptionCode <= _zz_statuses_0_exceptionCode_1;
        end
        if(_zz_123) begin
          statuses_6_exceptionCode <= _zz_statuses_0_exceptionCode_1;
        end
        if(_zz_124) begin
          statuses_7_exceptionCode <= _zz_statuses_0_exceptionCode_1;
        end
      end
      if(when_ReorderBuffer_l375_2) begin
        if(_zz_126) begin
          statuses_0_busy <= 1'b0;
        end
        if(_zz_127) begin
          statuses_1_busy <= 1'b0;
        end
        if(_zz_128) begin
          statuses_2_busy <= 1'b0;
        end
        if(_zz_129) begin
          statuses_3_busy <= 1'b0;
        end
        if(_zz_130) begin
          statuses_4_busy <= 1'b0;
        end
        if(_zz_131) begin
          statuses_5_busy <= 1'b0;
        end
        if(_zz_132) begin
          statuses_6_busy <= 1'b0;
        end
        if(_zz_133) begin
          statuses_7_busy <= 1'b0;
        end
        if(_zz_126) begin
          statuses_0_done <= 1'b1;
        end
        if(_zz_127) begin
          statuses_1_done <= 1'b1;
        end
        if(_zz_128) begin
          statuses_2_done <= 1'b1;
        end
        if(_zz_129) begin
          statuses_3_done <= 1'b1;
        end
        if(_zz_130) begin
          statuses_4_done <= 1'b1;
        end
        if(_zz_131) begin
          statuses_5_done <= 1'b1;
        end
        if(_zz_132) begin
          statuses_6_done <= 1'b1;
        end
        if(_zz_133) begin
          statuses_7_done <= 1'b1;
        end
        if(_zz_126) begin
          statuses_0_hasException <= io_writeback_2_exceptionOccurred;
        end
        if(_zz_127) begin
          statuses_1_hasException <= io_writeback_2_exceptionOccurred;
        end
        if(_zz_128) begin
          statuses_2_hasException <= io_writeback_2_exceptionOccurred;
        end
        if(_zz_129) begin
          statuses_3_hasException <= io_writeback_2_exceptionOccurred;
        end
        if(_zz_130) begin
          statuses_4_hasException <= io_writeback_2_exceptionOccurred;
        end
        if(_zz_131) begin
          statuses_5_hasException <= io_writeback_2_exceptionOccurred;
        end
        if(_zz_132) begin
          statuses_6_hasException <= io_writeback_2_exceptionOccurred;
        end
        if(_zz_133) begin
          statuses_7_hasException <= io_writeback_2_exceptionOccurred;
        end
        if(_zz_126) begin
          statuses_0_exceptionCode <= _zz_statuses_0_exceptionCode_2;
        end
        if(_zz_127) begin
          statuses_1_exceptionCode <= _zz_statuses_0_exceptionCode_2;
        end
        if(_zz_128) begin
          statuses_2_exceptionCode <= _zz_statuses_0_exceptionCode_2;
        end
        if(_zz_129) begin
          statuses_3_exceptionCode <= _zz_statuses_0_exceptionCode_2;
        end
        if(_zz_130) begin
          statuses_4_exceptionCode <= _zz_statuses_0_exceptionCode_2;
        end
        if(_zz_131) begin
          statuses_5_exceptionCode <= _zz_statuses_0_exceptionCode_2;
        end
        if(_zz_132) begin
          statuses_6_exceptionCode <= _zz_statuses_0_exceptionCode_2;
        end
        if(_zz_133) begin
          statuses_7_exceptionCode <= _zz_statuses_0_exceptionCode_2;
        end
      end
      if(when_ReorderBuffer_l375_3) begin
        if(_zz_135) begin
          statuses_0_busy <= 1'b0;
        end
        if(_zz_136) begin
          statuses_1_busy <= 1'b0;
        end
        if(_zz_137) begin
          statuses_2_busy <= 1'b0;
        end
        if(_zz_138) begin
          statuses_3_busy <= 1'b0;
        end
        if(_zz_139) begin
          statuses_4_busy <= 1'b0;
        end
        if(_zz_140) begin
          statuses_5_busy <= 1'b0;
        end
        if(_zz_141) begin
          statuses_6_busy <= 1'b0;
        end
        if(_zz_142) begin
          statuses_7_busy <= 1'b0;
        end
        if(_zz_135) begin
          statuses_0_done <= 1'b1;
        end
        if(_zz_136) begin
          statuses_1_done <= 1'b1;
        end
        if(_zz_137) begin
          statuses_2_done <= 1'b1;
        end
        if(_zz_138) begin
          statuses_3_done <= 1'b1;
        end
        if(_zz_139) begin
          statuses_4_done <= 1'b1;
        end
        if(_zz_140) begin
          statuses_5_done <= 1'b1;
        end
        if(_zz_141) begin
          statuses_6_done <= 1'b1;
        end
        if(_zz_142) begin
          statuses_7_done <= 1'b1;
        end
        if(_zz_135) begin
          statuses_0_hasException <= io_writeback_3_exceptionOccurred;
        end
        if(_zz_136) begin
          statuses_1_hasException <= io_writeback_3_exceptionOccurred;
        end
        if(_zz_137) begin
          statuses_2_hasException <= io_writeback_3_exceptionOccurred;
        end
        if(_zz_138) begin
          statuses_3_hasException <= io_writeback_3_exceptionOccurred;
        end
        if(_zz_139) begin
          statuses_4_hasException <= io_writeback_3_exceptionOccurred;
        end
        if(_zz_140) begin
          statuses_5_hasException <= io_writeback_3_exceptionOccurred;
        end
        if(_zz_141) begin
          statuses_6_hasException <= io_writeback_3_exceptionOccurred;
        end
        if(_zz_142) begin
          statuses_7_hasException <= io_writeback_3_exceptionOccurred;
        end
        if(_zz_135) begin
          statuses_0_exceptionCode <= _zz_statuses_0_exceptionCode_3;
        end
        if(_zz_136) begin
          statuses_1_exceptionCode <= _zz_statuses_0_exceptionCode_3;
        end
        if(_zz_137) begin
          statuses_2_exceptionCode <= _zz_statuses_0_exceptionCode_3;
        end
        if(_zz_138) begin
          statuses_3_exceptionCode <= _zz_statuses_0_exceptionCode_3;
        end
        if(_zz_139) begin
          statuses_4_exceptionCode <= _zz_statuses_0_exceptionCode_3;
        end
        if(_zz_140) begin
          statuses_5_exceptionCode <= _zz_statuses_0_exceptionCode_3;
        end
        if(_zz_141) begin
          statuses_6_exceptionCode <= _zz_statuses_0_exceptionCode_3;
        end
        if(_zz_142) begin
          statuses_7_exceptionCode <= _zz_statuses_0_exceptionCode_3;
        end
      end
      if(when_ReorderBuffer_l375_4) begin
        if(_zz_144) begin
          statuses_0_busy <= 1'b0;
        end
        if(_zz_145) begin
          statuses_1_busy <= 1'b0;
        end
        if(_zz_146) begin
          statuses_2_busy <= 1'b0;
        end
        if(_zz_147) begin
          statuses_3_busy <= 1'b0;
        end
        if(_zz_148) begin
          statuses_4_busy <= 1'b0;
        end
        if(_zz_149) begin
          statuses_5_busy <= 1'b0;
        end
        if(_zz_150) begin
          statuses_6_busy <= 1'b0;
        end
        if(_zz_151) begin
          statuses_7_busy <= 1'b0;
        end
        if(_zz_144) begin
          statuses_0_done <= 1'b1;
        end
        if(_zz_145) begin
          statuses_1_done <= 1'b1;
        end
        if(_zz_146) begin
          statuses_2_done <= 1'b1;
        end
        if(_zz_147) begin
          statuses_3_done <= 1'b1;
        end
        if(_zz_148) begin
          statuses_4_done <= 1'b1;
        end
        if(_zz_149) begin
          statuses_5_done <= 1'b1;
        end
        if(_zz_150) begin
          statuses_6_done <= 1'b1;
        end
        if(_zz_151) begin
          statuses_7_done <= 1'b1;
        end
        if(_zz_144) begin
          statuses_0_hasException <= io_writeback_4_exceptionOccurred;
        end
        if(_zz_145) begin
          statuses_1_hasException <= io_writeback_4_exceptionOccurred;
        end
        if(_zz_146) begin
          statuses_2_hasException <= io_writeback_4_exceptionOccurred;
        end
        if(_zz_147) begin
          statuses_3_hasException <= io_writeback_4_exceptionOccurred;
        end
        if(_zz_148) begin
          statuses_4_hasException <= io_writeback_4_exceptionOccurred;
        end
        if(_zz_149) begin
          statuses_5_hasException <= io_writeback_4_exceptionOccurred;
        end
        if(_zz_150) begin
          statuses_6_hasException <= io_writeback_4_exceptionOccurred;
        end
        if(_zz_151) begin
          statuses_7_hasException <= io_writeback_4_exceptionOccurred;
        end
        if(_zz_144) begin
          statuses_0_exceptionCode <= _zz_statuses_0_exceptionCode_4;
        end
        if(_zz_145) begin
          statuses_1_exceptionCode <= _zz_statuses_0_exceptionCode_4;
        end
        if(_zz_146) begin
          statuses_2_exceptionCode <= _zz_statuses_0_exceptionCode_4;
        end
        if(_zz_147) begin
          statuses_3_exceptionCode <= _zz_statuses_0_exceptionCode_4;
        end
        if(_zz_148) begin
          statuses_4_exceptionCode <= _zz_statuses_0_exceptionCode_4;
        end
        if(_zz_149) begin
          statuses_5_exceptionCode <= _zz_statuses_0_exceptionCode_4;
        end
        if(_zz_150) begin
          statuses_6_exceptionCode <= _zz_statuses_0_exceptionCode_4;
        end
        if(_zz_151) begin
          statuses_7_exceptionCode <= _zz_statuses_0_exceptionCode_4;
        end
      end
      if(io_flush_valid) begin
        case(io_flush_payload_reason)
          FlushReason_FULL_FLUSH : begin
            statuses_0_busy <= 1'b0;
            statuses_0_done <= 1'b0;
            statuses_0_hasException <= 1'b0;
            statuses_0_genBit <= 1'b0;
            statuses_1_busy <= 1'b0;
            statuses_1_done <= 1'b0;
            statuses_1_hasException <= 1'b0;
            statuses_1_genBit <= 1'b0;
            statuses_2_busy <= 1'b0;
            statuses_2_done <= 1'b0;
            statuses_2_hasException <= 1'b0;
            statuses_2_genBit <= 1'b0;
            statuses_3_busy <= 1'b0;
            statuses_3_done <= 1'b0;
            statuses_3_hasException <= 1'b0;
            statuses_3_genBit <= 1'b0;
            statuses_4_busy <= 1'b0;
            statuses_4_done <= 1'b0;
            statuses_4_hasException <= 1'b0;
            statuses_4_genBit <= 1'b0;
            statuses_5_busy <= 1'b0;
            statuses_5_done <= 1'b0;
            statuses_5_hasException <= 1'b0;
            statuses_5_genBit <= 1'b0;
            statuses_6_busy <= 1'b0;
            statuses_6_done <= 1'b0;
            statuses_6_hasException <= 1'b0;
            statuses_6_genBit <= 1'b0;
            statuses_7_busy <= 1'b0;
            statuses_7_done <= 1'b0;
            statuses_7_hasException <= 1'b0;
            statuses_7_genBit <= 1'b0;
          end
          FlushReason_ROLLBACK_TO_ROB_IDX : begin
            if(when_ReorderBuffer_l418) begin
              if(_zz_153) begin
                statuses_0_busy <= 1'b0;
              end
              if(_zz_154) begin
                statuses_1_busy <= 1'b0;
              end
              if(_zz_155) begin
                statuses_2_busy <= 1'b0;
              end
              if(_zz_156) begin
                statuses_3_busy <= 1'b0;
              end
              if(_zz_157) begin
                statuses_4_busy <= 1'b0;
              end
              if(_zz_158) begin
                statuses_5_busy <= 1'b0;
              end
              if(_zz_159) begin
                statuses_6_busy <= 1'b0;
              end
              if(_zz_160) begin
                statuses_7_busy <= 1'b0;
              end
              if(_zz_153) begin
                statuses_0_done <= 1'b0;
              end
              if(_zz_154) begin
                statuses_1_done <= 1'b0;
              end
              if(_zz_155) begin
                statuses_2_done <= 1'b0;
              end
              if(_zz_156) begin
                statuses_3_done <= 1'b0;
              end
              if(_zz_157) begin
                statuses_4_done <= 1'b0;
              end
              if(_zz_158) begin
                statuses_5_done <= 1'b0;
              end
              if(_zz_159) begin
                statuses_6_done <= 1'b0;
              end
              if(_zz_160) begin
                statuses_7_done <= 1'b0;
              end
              if(_zz_153) begin
                statuses_0_hasException <= 1'b0;
              end
              if(_zz_154) begin
                statuses_1_hasException <= 1'b0;
              end
              if(_zz_155) begin
                statuses_2_hasException <= 1'b0;
              end
              if(_zz_156) begin
                statuses_3_hasException <= 1'b0;
              end
              if(_zz_157) begin
                statuses_4_hasException <= 1'b0;
              end
              if(_zz_158) begin
                statuses_5_hasException <= 1'b0;
              end
              if(_zz_159) begin
                statuses_6_hasException <= 1'b0;
              end
              if(_zz_160) begin
                statuses_7_hasException <= 1'b0;
              end
            end
            if(when_ReorderBuffer_l418_1) begin
              if(_zz_162) begin
                statuses_0_busy <= 1'b0;
              end
              if(_zz_163) begin
                statuses_1_busy <= 1'b0;
              end
              if(_zz_164) begin
                statuses_2_busy <= 1'b0;
              end
              if(_zz_165) begin
                statuses_3_busy <= 1'b0;
              end
              if(_zz_166) begin
                statuses_4_busy <= 1'b0;
              end
              if(_zz_167) begin
                statuses_5_busy <= 1'b0;
              end
              if(_zz_168) begin
                statuses_6_busy <= 1'b0;
              end
              if(_zz_169) begin
                statuses_7_busy <= 1'b0;
              end
              if(_zz_162) begin
                statuses_0_done <= 1'b0;
              end
              if(_zz_163) begin
                statuses_1_done <= 1'b0;
              end
              if(_zz_164) begin
                statuses_2_done <= 1'b0;
              end
              if(_zz_165) begin
                statuses_3_done <= 1'b0;
              end
              if(_zz_166) begin
                statuses_4_done <= 1'b0;
              end
              if(_zz_167) begin
                statuses_5_done <= 1'b0;
              end
              if(_zz_168) begin
                statuses_6_done <= 1'b0;
              end
              if(_zz_169) begin
                statuses_7_done <= 1'b0;
              end
              if(_zz_162) begin
                statuses_0_hasException <= 1'b0;
              end
              if(_zz_163) begin
                statuses_1_hasException <= 1'b0;
              end
              if(_zz_164) begin
                statuses_2_hasException <= 1'b0;
              end
              if(_zz_165) begin
                statuses_3_hasException <= 1'b0;
              end
              if(_zz_166) begin
                statuses_4_hasException <= 1'b0;
              end
              if(_zz_167) begin
                statuses_5_hasException <= 1'b0;
              end
              if(_zz_168) begin
                statuses_6_hasException <= 1'b0;
              end
              if(_zz_169) begin
                statuses_7_hasException <= 1'b0;
              end
            end
            if(when_ReorderBuffer_l418_2) begin
              if(_zz_171) begin
                statuses_0_busy <= 1'b0;
              end
              if(_zz_172) begin
                statuses_1_busy <= 1'b0;
              end
              if(_zz_173) begin
                statuses_2_busy <= 1'b0;
              end
              if(_zz_174) begin
                statuses_3_busy <= 1'b0;
              end
              if(_zz_175) begin
                statuses_4_busy <= 1'b0;
              end
              if(_zz_176) begin
                statuses_5_busy <= 1'b0;
              end
              if(_zz_177) begin
                statuses_6_busy <= 1'b0;
              end
              if(_zz_178) begin
                statuses_7_busy <= 1'b0;
              end
              if(_zz_171) begin
                statuses_0_done <= 1'b0;
              end
              if(_zz_172) begin
                statuses_1_done <= 1'b0;
              end
              if(_zz_173) begin
                statuses_2_done <= 1'b0;
              end
              if(_zz_174) begin
                statuses_3_done <= 1'b0;
              end
              if(_zz_175) begin
                statuses_4_done <= 1'b0;
              end
              if(_zz_176) begin
                statuses_5_done <= 1'b0;
              end
              if(_zz_177) begin
                statuses_6_done <= 1'b0;
              end
              if(_zz_178) begin
                statuses_7_done <= 1'b0;
              end
              if(_zz_171) begin
                statuses_0_hasException <= 1'b0;
              end
              if(_zz_172) begin
                statuses_1_hasException <= 1'b0;
              end
              if(_zz_173) begin
                statuses_2_hasException <= 1'b0;
              end
              if(_zz_174) begin
                statuses_3_hasException <= 1'b0;
              end
              if(_zz_175) begin
                statuses_4_hasException <= 1'b0;
              end
              if(_zz_176) begin
                statuses_5_hasException <= 1'b0;
              end
              if(_zz_177) begin
                statuses_6_hasException <= 1'b0;
              end
              if(_zz_178) begin
                statuses_7_hasException <= 1'b0;
              end
            end
            if(when_ReorderBuffer_l418_3) begin
              if(_zz_180) begin
                statuses_0_busy <= 1'b0;
              end
              if(_zz_181) begin
                statuses_1_busy <= 1'b0;
              end
              if(_zz_182) begin
                statuses_2_busy <= 1'b0;
              end
              if(_zz_183) begin
                statuses_3_busy <= 1'b0;
              end
              if(_zz_184) begin
                statuses_4_busy <= 1'b0;
              end
              if(_zz_185) begin
                statuses_5_busy <= 1'b0;
              end
              if(_zz_186) begin
                statuses_6_busy <= 1'b0;
              end
              if(_zz_187) begin
                statuses_7_busy <= 1'b0;
              end
              if(_zz_180) begin
                statuses_0_done <= 1'b0;
              end
              if(_zz_181) begin
                statuses_1_done <= 1'b0;
              end
              if(_zz_182) begin
                statuses_2_done <= 1'b0;
              end
              if(_zz_183) begin
                statuses_3_done <= 1'b0;
              end
              if(_zz_184) begin
                statuses_4_done <= 1'b0;
              end
              if(_zz_185) begin
                statuses_5_done <= 1'b0;
              end
              if(_zz_186) begin
                statuses_6_done <= 1'b0;
              end
              if(_zz_187) begin
                statuses_7_done <= 1'b0;
              end
              if(_zz_180) begin
                statuses_0_hasException <= 1'b0;
              end
              if(_zz_181) begin
                statuses_1_hasException <= 1'b0;
              end
              if(_zz_182) begin
                statuses_2_hasException <= 1'b0;
              end
              if(_zz_183) begin
                statuses_3_hasException <= 1'b0;
              end
              if(_zz_184) begin
                statuses_4_hasException <= 1'b0;
              end
              if(_zz_185) begin
                statuses_5_hasException <= 1'b0;
              end
              if(_zz_186) begin
                statuses_6_hasException <= 1'b0;
              end
              if(_zz_187) begin
                statuses_7_hasException <= 1'b0;
              end
            end
            if(when_ReorderBuffer_l418_4) begin
              if(_zz_189) begin
                statuses_0_busy <= 1'b0;
              end
              if(_zz_190) begin
                statuses_1_busy <= 1'b0;
              end
              if(_zz_191) begin
                statuses_2_busy <= 1'b0;
              end
              if(_zz_192) begin
                statuses_3_busy <= 1'b0;
              end
              if(_zz_193) begin
                statuses_4_busy <= 1'b0;
              end
              if(_zz_194) begin
                statuses_5_busy <= 1'b0;
              end
              if(_zz_195) begin
                statuses_6_busy <= 1'b0;
              end
              if(_zz_196) begin
                statuses_7_busy <= 1'b0;
              end
              if(_zz_189) begin
                statuses_0_done <= 1'b0;
              end
              if(_zz_190) begin
                statuses_1_done <= 1'b0;
              end
              if(_zz_191) begin
                statuses_2_done <= 1'b0;
              end
              if(_zz_192) begin
                statuses_3_done <= 1'b0;
              end
              if(_zz_193) begin
                statuses_4_done <= 1'b0;
              end
              if(_zz_194) begin
                statuses_5_done <= 1'b0;
              end
              if(_zz_195) begin
                statuses_6_done <= 1'b0;
              end
              if(_zz_196) begin
                statuses_7_done <= 1'b0;
              end
              if(_zz_189) begin
                statuses_0_hasException <= 1'b0;
              end
              if(_zz_190) begin
                statuses_1_hasException <= 1'b0;
              end
              if(_zz_191) begin
                statuses_2_hasException <= 1'b0;
              end
              if(_zz_192) begin
                statuses_3_hasException <= 1'b0;
              end
              if(_zz_193) begin
                statuses_4_hasException <= 1'b0;
              end
              if(_zz_194) begin
                statuses_5_hasException <= 1'b0;
              end
              if(_zz_195) begin
                statuses_6_hasException <= 1'b0;
              end
              if(_zz_196) begin
                statuses_7_hasException <= 1'b0;
              end
            end
            if(when_ReorderBuffer_l418_5) begin
              if(_zz_198) begin
                statuses_0_busy <= 1'b0;
              end
              if(_zz_199) begin
                statuses_1_busy <= 1'b0;
              end
              if(_zz_200) begin
                statuses_2_busy <= 1'b0;
              end
              if(_zz_201) begin
                statuses_3_busy <= 1'b0;
              end
              if(_zz_202) begin
                statuses_4_busy <= 1'b0;
              end
              if(_zz_203) begin
                statuses_5_busy <= 1'b0;
              end
              if(_zz_204) begin
                statuses_6_busy <= 1'b0;
              end
              if(_zz_205) begin
                statuses_7_busy <= 1'b0;
              end
              if(_zz_198) begin
                statuses_0_done <= 1'b0;
              end
              if(_zz_199) begin
                statuses_1_done <= 1'b0;
              end
              if(_zz_200) begin
                statuses_2_done <= 1'b0;
              end
              if(_zz_201) begin
                statuses_3_done <= 1'b0;
              end
              if(_zz_202) begin
                statuses_4_done <= 1'b0;
              end
              if(_zz_203) begin
                statuses_5_done <= 1'b0;
              end
              if(_zz_204) begin
                statuses_6_done <= 1'b0;
              end
              if(_zz_205) begin
                statuses_7_done <= 1'b0;
              end
              if(_zz_198) begin
                statuses_0_hasException <= 1'b0;
              end
              if(_zz_199) begin
                statuses_1_hasException <= 1'b0;
              end
              if(_zz_200) begin
                statuses_2_hasException <= 1'b0;
              end
              if(_zz_201) begin
                statuses_3_hasException <= 1'b0;
              end
              if(_zz_202) begin
                statuses_4_hasException <= 1'b0;
              end
              if(_zz_203) begin
                statuses_5_hasException <= 1'b0;
              end
              if(_zz_204) begin
                statuses_6_hasException <= 1'b0;
              end
              if(_zz_205) begin
                statuses_7_hasException <= 1'b0;
              end
            end
            if(when_ReorderBuffer_l418_6) begin
              if(_zz_207) begin
                statuses_0_busy <= 1'b0;
              end
              if(_zz_208) begin
                statuses_1_busy <= 1'b0;
              end
              if(_zz_209) begin
                statuses_2_busy <= 1'b0;
              end
              if(_zz_210) begin
                statuses_3_busy <= 1'b0;
              end
              if(_zz_211) begin
                statuses_4_busy <= 1'b0;
              end
              if(_zz_212) begin
                statuses_5_busy <= 1'b0;
              end
              if(_zz_213) begin
                statuses_6_busy <= 1'b0;
              end
              if(_zz_214) begin
                statuses_7_busy <= 1'b0;
              end
              if(_zz_207) begin
                statuses_0_done <= 1'b0;
              end
              if(_zz_208) begin
                statuses_1_done <= 1'b0;
              end
              if(_zz_209) begin
                statuses_2_done <= 1'b0;
              end
              if(_zz_210) begin
                statuses_3_done <= 1'b0;
              end
              if(_zz_211) begin
                statuses_4_done <= 1'b0;
              end
              if(_zz_212) begin
                statuses_5_done <= 1'b0;
              end
              if(_zz_213) begin
                statuses_6_done <= 1'b0;
              end
              if(_zz_214) begin
                statuses_7_done <= 1'b0;
              end
              if(_zz_207) begin
                statuses_0_hasException <= 1'b0;
              end
              if(_zz_208) begin
                statuses_1_hasException <= 1'b0;
              end
              if(_zz_209) begin
                statuses_2_hasException <= 1'b0;
              end
              if(_zz_210) begin
                statuses_3_hasException <= 1'b0;
              end
              if(_zz_211) begin
                statuses_4_hasException <= 1'b0;
              end
              if(_zz_212) begin
                statuses_5_hasException <= 1'b0;
              end
              if(_zz_213) begin
                statuses_6_hasException <= 1'b0;
              end
              if(_zz_214) begin
                statuses_7_hasException <= 1'b0;
              end
            end
            if(when_ReorderBuffer_l418_7) begin
              if(_zz_216) begin
                statuses_0_busy <= 1'b0;
              end
              if(_zz_217) begin
                statuses_1_busy <= 1'b0;
              end
              if(_zz_218) begin
                statuses_2_busy <= 1'b0;
              end
              if(_zz_219) begin
                statuses_3_busy <= 1'b0;
              end
              if(_zz_220) begin
                statuses_4_busy <= 1'b0;
              end
              if(_zz_221) begin
                statuses_5_busy <= 1'b0;
              end
              if(_zz_222) begin
                statuses_6_busy <= 1'b0;
              end
              if(_zz_223) begin
                statuses_7_busy <= 1'b0;
              end
              if(_zz_216) begin
                statuses_0_done <= 1'b0;
              end
              if(_zz_217) begin
                statuses_1_done <= 1'b0;
              end
              if(_zz_218) begin
                statuses_2_done <= 1'b0;
              end
              if(_zz_219) begin
                statuses_3_done <= 1'b0;
              end
              if(_zz_220) begin
                statuses_4_done <= 1'b0;
              end
              if(_zz_221) begin
                statuses_5_done <= 1'b0;
              end
              if(_zz_222) begin
                statuses_6_done <= 1'b0;
              end
              if(_zz_223) begin
                statuses_7_done <= 1'b0;
              end
              if(_zz_216) begin
                statuses_0_hasException <= 1'b0;
              end
              if(_zz_217) begin
                statuses_1_hasException <= 1'b0;
              end
              if(_zz_218) begin
                statuses_2_hasException <= 1'b0;
              end
              if(_zz_219) begin
                statuses_3_hasException <= 1'b0;
              end
              if(_zz_220) begin
                statuses_4_hasException <= 1'b0;
              end
              if(_zz_221) begin
                statuses_5_hasException <= 1'b0;
              end
              if(_zz_222) begin
                statuses_6_hasException <= 1'b0;
              end
              if(_zz_223) begin
                statuses_7_hasException <= 1'b0;
              end
            end
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(posedge clk) begin
    if(when_ReorderBuffer_l375) begin
      if(_zz_108) begin
        statuses_0_isMispredictedBranch <= io_writeback_0_isMispredictedBranch;
      end
      if(_zz_109) begin
        statuses_1_isMispredictedBranch <= io_writeback_0_isMispredictedBranch;
      end
      if(_zz_110) begin
        statuses_2_isMispredictedBranch <= io_writeback_0_isMispredictedBranch;
      end
      if(_zz_111) begin
        statuses_3_isMispredictedBranch <= io_writeback_0_isMispredictedBranch;
      end
      if(_zz_112) begin
        statuses_4_isMispredictedBranch <= io_writeback_0_isMispredictedBranch;
      end
      if(_zz_113) begin
        statuses_5_isMispredictedBranch <= io_writeback_0_isMispredictedBranch;
      end
      if(_zz_114) begin
        statuses_6_isMispredictedBranch <= io_writeback_0_isMispredictedBranch;
      end
      if(_zz_115) begin
        statuses_7_isMispredictedBranch <= io_writeback_0_isMispredictedBranch;
      end
      if(_zz_108) begin
        statuses_0_isTaken <= io_writeback_0_isTaken;
      end
      if(_zz_109) begin
        statuses_1_isTaken <= io_writeback_0_isTaken;
      end
      if(_zz_110) begin
        statuses_2_isTaken <= io_writeback_0_isTaken;
      end
      if(_zz_111) begin
        statuses_3_isTaken <= io_writeback_0_isTaken;
      end
      if(_zz_112) begin
        statuses_4_isTaken <= io_writeback_0_isTaken;
      end
      if(_zz_113) begin
        statuses_5_isTaken <= io_writeback_0_isTaken;
      end
      if(_zz_114) begin
        statuses_6_isTaken <= io_writeback_0_isTaken;
      end
      if(_zz_115) begin
        statuses_7_isTaken <= io_writeback_0_isTaken;
      end
      if(_zz_108) begin
        statuses_0_result <= io_writeback_0_result;
      end
      if(_zz_109) begin
        statuses_1_result <= io_writeback_0_result;
      end
      if(_zz_110) begin
        statuses_2_result <= io_writeback_0_result;
      end
      if(_zz_111) begin
        statuses_3_result <= io_writeback_0_result;
      end
      if(_zz_112) begin
        statuses_4_result <= io_writeback_0_result;
      end
      if(_zz_113) begin
        statuses_5_result <= io_writeback_0_result;
      end
      if(_zz_114) begin
        statuses_6_result <= io_writeback_0_result;
      end
      if(_zz_115) begin
        statuses_7_result <= io_writeback_0_result;
      end
    end
    if(when_ReorderBuffer_l375_1) begin
      if(_zz_117) begin
        statuses_0_isMispredictedBranch <= io_writeback_1_isMispredictedBranch;
      end
      if(_zz_118) begin
        statuses_1_isMispredictedBranch <= io_writeback_1_isMispredictedBranch;
      end
      if(_zz_119) begin
        statuses_2_isMispredictedBranch <= io_writeback_1_isMispredictedBranch;
      end
      if(_zz_120) begin
        statuses_3_isMispredictedBranch <= io_writeback_1_isMispredictedBranch;
      end
      if(_zz_121) begin
        statuses_4_isMispredictedBranch <= io_writeback_1_isMispredictedBranch;
      end
      if(_zz_122) begin
        statuses_5_isMispredictedBranch <= io_writeback_1_isMispredictedBranch;
      end
      if(_zz_123) begin
        statuses_6_isMispredictedBranch <= io_writeback_1_isMispredictedBranch;
      end
      if(_zz_124) begin
        statuses_7_isMispredictedBranch <= io_writeback_1_isMispredictedBranch;
      end
      if(_zz_117) begin
        statuses_0_isTaken <= io_writeback_1_isTaken;
      end
      if(_zz_118) begin
        statuses_1_isTaken <= io_writeback_1_isTaken;
      end
      if(_zz_119) begin
        statuses_2_isTaken <= io_writeback_1_isTaken;
      end
      if(_zz_120) begin
        statuses_3_isTaken <= io_writeback_1_isTaken;
      end
      if(_zz_121) begin
        statuses_4_isTaken <= io_writeback_1_isTaken;
      end
      if(_zz_122) begin
        statuses_5_isTaken <= io_writeback_1_isTaken;
      end
      if(_zz_123) begin
        statuses_6_isTaken <= io_writeback_1_isTaken;
      end
      if(_zz_124) begin
        statuses_7_isTaken <= io_writeback_1_isTaken;
      end
      if(_zz_117) begin
        statuses_0_result <= io_writeback_1_result;
      end
      if(_zz_118) begin
        statuses_1_result <= io_writeback_1_result;
      end
      if(_zz_119) begin
        statuses_2_result <= io_writeback_1_result;
      end
      if(_zz_120) begin
        statuses_3_result <= io_writeback_1_result;
      end
      if(_zz_121) begin
        statuses_4_result <= io_writeback_1_result;
      end
      if(_zz_122) begin
        statuses_5_result <= io_writeback_1_result;
      end
      if(_zz_123) begin
        statuses_6_result <= io_writeback_1_result;
      end
      if(_zz_124) begin
        statuses_7_result <= io_writeback_1_result;
      end
    end
    if(when_ReorderBuffer_l375_2) begin
      if(_zz_126) begin
        statuses_0_isMispredictedBranch <= io_writeback_2_isMispredictedBranch;
      end
      if(_zz_127) begin
        statuses_1_isMispredictedBranch <= io_writeback_2_isMispredictedBranch;
      end
      if(_zz_128) begin
        statuses_2_isMispredictedBranch <= io_writeback_2_isMispredictedBranch;
      end
      if(_zz_129) begin
        statuses_3_isMispredictedBranch <= io_writeback_2_isMispredictedBranch;
      end
      if(_zz_130) begin
        statuses_4_isMispredictedBranch <= io_writeback_2_isMispredictedBranch;
      end
      if(_zz_131) begin
        statuses_5_isMispredictedBranch <= io_writeback_2_isMispredictedBranch;
      end
      if(_zz_132) begin
        statuses_6_isMispredictedBranch <= io_writeback_2_isMispredictedBranch;
      end
      if(_zz_133) begin
        statuses_7_isMispredictedBranch <= io_writeback_2_isMispredictedBranch;
      end
      if(_zz_126) begin
        statuses_0_isTaken <= io_writeback_2_isTaken;
      end
      if(_zz_127) begin
        statuses_1_isTaken <= io_writeback_2_isTaken;
      end
      if(_zz_128) begin
        statuses_2_isTaken <= io_writeback_2_isTaken;
      end
      if(_zz_129) begin
        statuses_3_isTaken <= io_writeback_2_isTaken;
      end
      if(_zz_130) begin
        statuses_4_isTaken <= io_writeback_2_isTaken;
      end
      if(_zz_131) begin
        statuses_5_isTaken <= io_writeback_2_isTaken;
      end
      if(_zz_132) begin
        statuses_6_isTaken <= io_writeback_2_isTaken;
      end
      if(_zz_133) begin
        statuses_7_isTaken <= io_writeback_2_isTaken;
      end
      if(_zz_126) begin
        statuses_0_result <= io_writeback_2_result;
      end
      if(_zz_127) begin
        statuses_1_result <= io_writeback_2_result;
      end
      if(_zz_128) begin
        statuses_2_result <= io_writeback_2_result;
      end
      if(_zz_129) begin
        statuses_3_result <= io_writeback_2_result;
      end
      if(_zz_130) begin
        statuses_4_result <= io_writeback_2_result;
      end
      if(_zz_131) begin
        statuses_5_result <= io_writeback_2_result;
      end
      if(_zz_132) begin
        statuses_6_result <= io_writeback_2_result;
      end
      if(_zz_133) begin
        statuses_7_result <= io_writeback_2_result;
      end
    end
    if(when_ReorderBuffer_l375_3) begin
      if(_zz_135) begin
        statuses_0_isMispredictedBranch <= io_writeback_3_isMispredictedBranch;
      end
      if(_zz_136) begin
        statuses_1_isMispredictedBranch <= io_writeback_3_isMispredictedBranch;
      end
      if(_zz_137) begin
        statuses_2_isMispredictedBranch <= io_writeback_3_isMispredictedBranch;
      end
      if(_zz_138) begin
        statuses_3_isMispredictedBranch <= io_writeback_3_isMispredictedBranch;
      end
      if(_zz_139) begin
        statuses_4_isMispredictedBranch <= io_writeback_3_isMispredictedBranch;
      end
      if(_zz_140) begin
        statuses_5_isMispredictedBranch <= io_writeback_3_isMispredictedBranch;
      end
      if(_zz_141) begin
        statuses_6_isMispredictedBranch <= io_writeback_3_isMispredictedBranch;
      end
      if(_zz_142) begin
        statuses_7_isMispredictedBranch <= io_writeback_3_isMispredictedBranch;
      end
      if(_zz_135) begin
        statuses_0_isTaken <= io_writeback_3_isTaken;
      end
      if(_zz_136) begin
        statuses_1_isTaken <= io_writeback_3_isTaken;
      end
      if(_zz_137) begin
        statuses_2_isTaken <= io_writeback_3_isTaken;
      end
      if(_zz_138) begin
        statuses_3_isTaken <= io_writeback_3_isTaken;
      end
      if(_zz_139) begin
        statuses_4_isTaken <= io_writeback_3_isTaken;
      end
      if(_zz_140) begin
        statuses_5_isTaken <= io_writeback_3_isTaken;
      end
      if(_zz_141) begin
        statuses_6_isTaken <= io_writeback_3_isTaken;
      end
      if(_zz_142) begin
        statuses_7_isTaken <= io_writeback_3_isTaken;
      end
      if(_zz_135) begin
        statuses_0_result <= io_writeback_3_result;
      end
      if(_zz_136) begin
        statuses_1_result <= io_writeback_3_result;
      end
      if(_zz_137) begin
        statuses_2_result <= io_writeback_3_result;
      end
      if(_zz_138) begin
        statuses_3_result <= io_writeback_3_result;
      end
      if(_zz_139) begin
        statuses_4_result <= io_writeback_3_result;
      end
      if(_zz_140) begin
        statuses_5_result <= io_writeback_3_result;
      end
      if(_zz_141) begin
        statuses_6_result <= io_writeback_3_result;
      end
      if(_zz_142) begin
        statuses_7_result <= io_writeback_3_result;
      end
    end
    if(when_ReorderBuffer_l375_4) begin
      if(_zz_144) begin
        statuses_0_isMispredictedBranch <= io_writeback_4_isMispredictedBranch;
      end
      if(_zz_145) begin
        statuses_1_isMispredictedBranch <= io_writeback_4_isMispredictedBranch;
      end
      if(_zz_146) begin
        statuses_2_isMispredictedBranch <= io_writeback_4_isMispredictedBranch;
      end
      if(_zz_147) begin
        statuses_3_isMispredictedBranch <= io_writeback_4_isMispredictedBranch;
      end
      if(_zz_148) begin
        statuses_4_isMispredictedBranch <= io_writeback_4_isMispredictedBranch;
      end
      if(_zz_149) begin
        statuses_5_isMispredictedBranch <= io_writeback_4_isMispredictedBranch;
      end
      if(_zz_150) begin
        statuses_6_isMispredictedBranch <= io_writeback_4_isMispredictedBranch;
      end
      if(_zz_151) begin
        statuses_7_isMispredictedBranch <= io_writeback_4_isMispredictedBranch;
      end
      if(_zz_144) begin
        statuses_0_isTaken <= io_writeback_4_isTaken;
      end
      if(_zz_145) begin
        statuses_1_isTaken <= io_writeback_4_isTaken;
      end
      if(_zz_146) begin
        statuses_2_isTaken <= io_writeback_4_isTaken;
      end
      if(_zz_147) begin
        statuses_3_isTaken <= io_writeback_4_isTaken;
      end
      if(_zz_148) begin
        statuses_4_isTaken <= io_writeback_4_isTaken;
      end
      if(_zz_149) begin
        statuses_5_isTaken <= io_writeback_4_isTaken;
      end
      if(_zz_150) begin
        statuses_6_isTaken <= io_writeback_4_isTaken;
      end
      if(_zz_151) begin
        statuses_7_isTaken <= io_writeback_4_isTaken;
      end
      if(_zz_144) begin
        statuses_0_result <= io_writeback_4_result;
      end
      if(_zz_145) begin
        statuses_1_result <= io_writeback_4_result;
      end
      if(_zz_146) begin
        statuses_2_result <= io_writeback_4_result;
      end
      if(_zz_147) begin
        statuses_3_result <= io_writeback_4_result;
      end
      if(_zz_148) begin
        statuses_4_result <= io_writeback_4_result;
      end
      if(_zz_149) begin
        statuses_5_result <= io_writeback_4_result;
      end
      if(_zz_150) begin
        statuses_6_result <= io_writeback_4_result;
      end
      if(_zz_151) begin
        statuses_7_result <= io_writeback_4_result;
      end
    end
  end


endmodule

module StreamFifo_11 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_pc,
  input  wire [31:0]   io_push_payload_instruction,
  input  wire          io_push_payload_predecode_isBranch,
  input  wire          io_push_payload_predecode_isJump,
  input  wire          io_push_payload_predecode_isDirectJump,
  input  wire [31:0]   io_push_payload_predecode_jumpOffset,
  input  wire          io_push_payload_predecode_isIdle,
  input  wire          io_push_payload_bpuPrediction_isTaken,
  input  wire [31:0]   io_push_payload_bpuPrediction_target,
  input  wire          io_push_payload_bpuPrediction_wasPredicted,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_pc,
  output wire [31:0]   io_pop_payload_instruction,
  output wire          io_pop_payload_predecode_isBranch,
  output wire          io_pop_payload_predecode_isJump,
  output wire          io_pop_payload_predecode_isDirectJump,
  output wire [31:0]   io_pop_payload_predecode_jumpOffset,
  output wire          io_pop_payload_predecode_isIdle,
  output wire          io_pop_payload_bpuPrediction_isTaken,
  output wire [31:0]   io_pop_payload_bpuPrediction_target,
  output wire          io_pop_payload_bpuPrediction_wasPredicted,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [133:0]  logic_ram_spinal_port1;
  wire       [133:0]  _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1455;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [1:0]    logic_push_onRam_write_payload_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_pc;
  wire       [31:0]   logic_push_onRam_write_payload_data_instruction;
  wire                logic_push_onRam_write_payload_data_predecode_isBranch;
  wire                logic_push_onRam_write_payload_data_predecode_isJump;
  wire                logic_push_onRam_write_payload_data_predecode_isDirectJump;
  wire       [31:0]   logic_push_onRam_write_payload_data_predecode_jumpOffset;
  wire                logic_push_onRam_write_payload_data_predecode_isIdle;
  wire                logic_push_onRam_write_payload_data_bpuPrediction_isTaken;
  wire       [31:0]   logic_push_onRam_write_payload_data_bpuPrediction_target;
  wire                logic_push_onRam_write_payload_data_bpuPrediction_wasPredicted;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [1:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [1:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [1:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l477;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [1:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [31:0]   logic_pop_sync_readPort_rsp_pc;
  wire       [31:0]   logic_pop_sync_readPort_rsp_instruction;
  wire                logic_pop_sync_readPort_rsp_predecode_isBranch;
  wire                logic_pop_sync_readPort_rsp_predecode_isJump;
  wire                logic_pop_sync_readPort_rsp_predecode_isDirectJump;
  wire       [31:0]   logic_pop_sync_readPort_rsp_predecode_jumpOffset;
  wire                logic_pop_sync_readPort_rsp_predecode_isIdle;
  wire                logic_pop_sync_readPort_rsp_bpuPrediction_isTaken;
  wire       [31:0]   logic_pop_sync_readPort_rsp_bpuPrediction_target;
  wire                logic_pop_sync_readPort_rsp_bpuPrediction_wasPredicted;
  wire       [133:0]  _zz_logic_pop_sync_readPort_rsp_pc;
  wire       [35:0]   _zz_logic_pop_sync_readPort_rsp_predecode_isBranch;
  wire       [33:0]   _zz_logic_pop_sync_readPort_rsp_bpuPrediction_isTaken;
  wire                logic_pop_addressGen_toFlowFire_valid;
  wire       [1:0]    logic_pop_addressGen_toFlowFire_payload;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_pc;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_instruction;
  wire                logic_pop_sync_readArbitation_translated_payload_predecode_isBranch;
  wire                logic_pop_sync_readArbitation_translated_payload_predecode_isJump;
  wire                logic_pop_sync_readArbitation_translated_payload_predecode_isDirectJump;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_predecode_jumpOffset;
  wire                logic_pop_sync_readArbitation_translated_payload_predecode_isIdle;
  wire                logic_pop_sync_readArbitation_translated_payload_bpuPrediction_isTaken;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_bpuPrediction_target;
  wire                logic_pop_sync_readArbitation_translated_payload_bpuPrediction_wasPredicted;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [2:0]    logic_pop_sync_popReg;
  (* ram_style = "block" *) reg [133:0] logic_ram [0:3];

  assign _zz_logic_ram_port = {{logic_push_onRam_write_payload_data_bpuPrediction_wasPredicted,{logic_push_onRam_write_payload_data_bpuPrediction_target,logic_push_onRam_write_payload_data_bpuPrediction_isTaken}},{{logic_push_onRam_write_payload_data_predecode_isIdle,{logic_push_onRam_write_payload_data_predecode_jumpOffset,{logic_push_onRam_write_payload_data_predecode_isDirectJump,{logic_push_onRam_write_payload_data_predecode_isJump,logic_push_onRam_write_payload_data_predecode_isBranch}}}},{logic_push_onRam_write_payload_data_instruction,logic_push_onRam_write_payload_data_pc}}};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1455 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 3'b100) == 3'b000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[1:0];
  assign logic_push_onRam_write_payload_data_pc = io_push_payload_pc;
  assign logic_push_onRam_write_payload_data_instruction = io_push_payload_instruction;
  assign logic_push_onRam_write_payload_data_predecode_isBranch = io_push_payload_predecode_isBranch;
  assign logic_push_onRam_write_payload_data_predecode_isJump = io_push_payload_predecode_isJump;
  assign logic_push_onRam_write_payload_data_predecode_isDirectJump = io_push_payload_predecode_isDirectJump;
  assign logic_push_onRam_write_payload_data_predecode_jumpOffset = io_push_payload_predecode_jumpOffset;
  assign logic_push_onRam_write_payload_data_predecode_isIdle = io_push_payload_predecode_isIdle;
  assign logic_push_onRam_write_payload_data_bpuPrediction_isTaken = io_push_payload_bpuPrediction_isTaken;
  assign logic_push_onRam_write_payload_data_bpuPrediction_target = io_push_payload_bpuPrediction_target;
  assign logic_push_onRam_write_payload_data_bpuPrediction_wasPredicted = io_push_payload_bpuPrediction_wasPredicted;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[1:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l477) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_pc = logic_ram_spinal_port1;
  assign _zz_logic_pop_sync_readPort_rsp_predecode_isBranch = _zz_logic_pop_sync_readPort_rsp_pc[99 : 64];
  assign _zz_logic_pop_sync_readPort_rsp_bpuPrediction_isTaken = _zz_logic_pop_sync_readPort_rsp_pc[133 : 100];
  assign logic_pop_sync_readPort_rsp_pc = _zz_logic_pop_sync_readPort_rsp_pc[31 : 0];
  assign logic_pop_sync_readPort_rsp_instruction = _zz_logic_pop_sync_readPort_rsp_pc[63 : 32];
  assign logic_pop_sync_readPort_rsp_predecode_isBranch = _zz_logic_pop_sync_readPort_rsp_predecode_isBranch[0];
  assign logic_pop_sync_readPort_rsp_predecode_isJump = _zz_logic_pop_sync_readPort_rsp_predecode_isBranch[1];
  assign logic_pop_sync_readPort_rsp_predecode_isDirectJump = _zz_logic_pop_sync_readPort_rsp_predecode_isBranch[2];
  assign logic_pop_sync_readPort_rsp_predecode_jumpOffset = _zz_logic_pop_sync_readPort_rsp_predecode_isBranch[34 : 3];
  assign logic_pop_sync_readPort_rsp_predecode_isIdle = _zz_logic_pop_sync_readPort_rsp_predecode_isBranch[35];
  assign logic_pop_sync_readPort_rsp_bpuPrediction_isTaken = _zz_logic_pop_sync_readPort_rsp_bpuPrediction_isTaken[0];
  assign logic_pop_sync_readPort_rsp_bpuPrediction_target = _zz_logic_pop_sync_readPort_rsp_bpuPrediction_isTaken[32 : 1];
  assign logic_pop_sync_readPort_rsp_bpuPrediction_wasPredicted = _zz_logic_pop_sync_readPort_rsp_bpuPrediction_isTaken[33];
  assign logic_pop_addressGen_toFlowFire_valid = logic_pop_addressGen_fire;
  assign logic_pop_addressGen_toFlowFire_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_toFlowFire_valid;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_toFlowFire_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_pc = logic_pop_sync_readPort_rsp_pc;
  assign logic_pop_sync_readArbitation_translated_payload_instruction = logic_pop_sync_readPort_rsp_instruction;
  assign logic_pop_sync_readArbitation_translated_payload_predecode_isBranch = logic_pop_sync_readPort_rsp_predecode_isBranch;
  assign logic_pop_sync_readArbitation_translated_payload_predecode_isJump = logic_pop_sync_readPort_rsp_predecode_isJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecode_isDirectJump = logic_pop_sync_readPort_rsp_predecode_isDirectJump;
  assign logic_pop_sync_readArbitation_translated_payload_predecode_jumpOffset = logic_pop_sync_readPort_rsp_predecode_jumpOffset;
  assign logic_pop_sync_readArbitation_translated_payload_predecode_isIdle = logic_pop_sync_readPort_rsp_predecode_isIdle;
  assign logic_pop_sync_readArbitation_translated_payload_bpuPrediction_isTaken = logic_pop_sync_readPort_rsp_bpuPrediction_isTaken;
  assign logic_pop_sync_readArbitation_translated_payload_bpuPrediction_target = logic_pop_sync_readPort_rsp_bpuPrediction_target;
  assign logic_pop_sync_readArbitation_translated_payload_bpuPrediction_wasPredicted = logic_pop_sync_readPort_rsp_bpuPrediction_wasPredicted;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_pc = logic_pop_sync_readArbitation_translated_payload_pc;
  assign io_pop_payload_instruction = logic_pop_sync_readArbitation_translated_payload_instruction;
  assign io_pop_payload_predecode_isBranch = logic_pop_sync_readArbitation_translated_payload_predecode_isBranch;
  assign io_pop_payload_predecode_isJump = logic_pop_sync_readArbitation_translated_payload_predecode_isJump;
  assign io_pop_payload_predecode_isDirectJump = logic_pop_sync_readArbitation_translated_payload_predecode_isDirectJump;
  assign io_pop_payload_predecode_jumpOffset = logic_pop_sync_readArbitation_translated_payload_predecode_jumpOffset;
  assign io_pop_payload_predecode_isIdle = logic_pop_sync_readArbitation_translated_payload_predecode_isIdle;
  assign io_pop_payload_bpuPrediction_isTaken = logic_pop_sync_readArbitation_translated_payload_bpuPrediction_isTaken;
  assign io_pop_payload_bpuPrediction_target = logic_pop_sync_readArbitation_translated_payload_bpuPrediction_target;
  assign io_pop_payload_bpuPrediction_wasPredicted = logic_pop_sync_readArbitation_translated_payload_bpuPrediction_wasPredicted;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b100 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 3'b000;
    end else begin
      if(when_Stream_l1455) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 3'b000;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module OneShot (
  input  wire          io_triggerIn,
  output reg           io_pulseOut,
  input  wire          clk,
  input  wire          reset
);

  reg                 hasFired;
  wire                when_Debug_l150;

  always @(*) begin
    io_pulseOut = 1'b0;
    if(when_Debug_l150) begin
      io_pulseOut = 1'b1;
    end
  end

  assign when_Debug_l150 = (io_triggerIn && (! hasFired));
  always @(posedge clk) begin
    if(reset) begin
      hasFired <= 1'b0;
    end else begin
      if(when_Debug_l150) begin
        hasFired <= 1'b1;
      end
    end
  end


endmodule

module DataCache (
  input  wire          io_load_cmd_valid,
  output wire          io_load_cmd_ready,
  input  wire [31:0]   io_load_cmd_payload_virtual,
  input  wire [1:0]    io_load_cmd_payload_size,
  input  wire          io_load_cmd_payload_redoOnDataHazard,
  input  wire [2:0]    io_load_cmd_payload_transactionId,
  input  wire [2:0]    io_load_cmd_payload_id,
  input  wire [31:0]   io_load_translated_physical,
  input  wire          io_load_translated_abord,
  input  wire [2:0]    io_load_cancels,
  output wire          io_load_rsp_valid,
  output wire [31:0]   io_load_rsp_payload_data,
  output wire          io_load_rsp_payload_fault,
  output wire          io_load_rsp_payload_redo,
  output wire [7:0]    io_load_rsp_payload_refillSlot,
  output wire          io_load_rsp_payload_refillSlotAny,
  output wire [2:0]    io_load_rsp_payload_id,
  input  wire          io_store_cmd_valid,
  output wire          io_store_cmd_ready,
  input  wire [31:0]   io_store_cmd_payload_address,
  input  wire [31:0]   io_store_cmd_payload_data,
  input  wire [3:0]    io_store_cmd_payload_mask,
  input  wire          io_store_cmd_payload_io,
  input  wire          io_store_cmd_payload_flush,
  input  wire          io_store_cmd_payload_flushFree,
  input  wire          io_store_cmd_payload_prefetch,
  input  wire [2:0]    io_store_cmd_payload_id,
  output wire          io_store_rsp_valid,
  output wire          io_store_rsp_payload_fault,
  output wire          io_store_rsp_payload_redo,
  output wire [7:0]    io_store_rsp_payload_refillSlot,
  output wire          io_store_rsp_payload_refillSlotAny,
  output wire          io_store_rsp_payload_flush,
  output wire          io_store_rsp_payload_prefetch,
  output wire [31:0]   io_store_rsp_payload_address,
  output wire          io_store_rsp_payload_io,
  output wire [2:0]    io_store_rsp_payload_id,
  output wire          io_mem_read_cmd_valid,
  input  wire          io_mem_read_cmd_ready,
  output wire [2:0]    io_mem_read_cmd_payload_id,
  output wire [31:0]   io_mem_read_cmd_payload_address,
  input  wire          io_mem_read_rsp_valid,
  output wire          io_mem_read_rsp_ready,
  input  wire [2:0]    io_mem_read_rsp_payload_id,
  input  wire [31:0]   io_mem_read_rsp_payload_data,
  input  wire          io_mem_read_rsp_payload_error,
  output wire          io_mem_write_cmd_valid,
  input  wire          io_mem_write_cmd_ready,
  output wire          io_mem_write_cmd_payload_last,
  output wire [31:0]   io_mem_write_cmd_payload_fragment_address,
  output wire [31:0]   io_mem_write_cmd_payload_fragment_data,
  output wire [2:0]    io_mem_write_cmd_payload_fragment_id,
  input  wire          io_mem_write_rsp_valid,
  input  wire          io_mem_write_rsp_payload_error,
  input  wire [2:0]    io_mem_write_rsp_payload_id,
  output reg  [7:0]    io_refillCompletions,
  output wire          io_refillEvent,
  output wire          io_writebackEvent,
  output wire          io_writebackBusy,
  input  wire          clk,
  input  wire          reset
);

  reg        [31:0]   banks_0_mem_spinal_port1;
  reg        [31:0]   banks_1_mem_spinal_port1;
  wire       [24:0]   ways_0_mem_spinal_port1;
  wire       [24:0]   ways_0_mem_spinal_port2;
  wire       [24:0]   ways_1_mem_spinal_port1;
  wire       [24:0]   ways_1_mem_spinal_port2;
  wire       [1:0]    status_mem_spinal_port1;
  wire       [1:0]    status_mem_spinal_port2;
  reg        [31:0]   writeback_victimBuffer_spinal_port1;
  wire       [24:0]   _zz_ways_0_mem_port;
  wire                _zz_ways_0_mem_port_1;
  wire       [24:0]   _zz_ways_1_mem_port;
  wire                _zz_ways_1_mem_port_1;
  wire       [1:0]    _zz_status_mem_port;
  wire       [0:0]    _zz_status_loadRead_rsp_0_dirty_1;
  wire       [0:0]    _zz_status_loadRead_rsp_1_dirty;
  wire       [0:0]    _zz_status_storeRead_rsp_0_dirty_1;
  wire       [0:0]    _zz_status_storeRead_rsp_1_dirty;
  wire       [7:0]    _zz__zz_refill_free_1;
  wire                _zz_refill_read_arbiter_oh;
  wire       [0:0]    _zz_refill_read_arbiter_oh_1;
  wire       [4:0]    _zz_refill_read_arbiter_oh_2;
  wire                _zz_refill_read_arbiter_oh_3;
  wire       [0:0]    _zz_refill_read_arbiter_oh_4;
  wire       [2:0]    _zz_refill_read_arbiter_oh_5;
  wire                _zz_refill_read_arbiter_oh_6;
  wire       [0:0]    _zz_refill_read_arbiter_oh_7;
  wire       [0:0]    _zz_refill_read_arbiter_oh_8;
  wire       [0:0]    _zz_refill_read_arbiter_oh_9;
  wire       [5:0]    _zz_refill_read_arbiter_oh_10;
  wire                _zz_refill_read_arbiter_oh_11;
  wire       [0:0]    _zz_refill_read_arbiter_oh_12;
  wire       [3:0]    _zz_refill_read_arbiter_oh_13;
  wire                _zz_refill_read_arbiter_oh_14;
  wire       [0:0]    _zz_refill_read_arbiter_oh_15;
  wire       [1:0]    _zz_refill_read_arbiter_oh_16;
  wire                _zz_refill_read_arbiter_oh_17;
  wire                _zz_refill_read_arbiter_oh_18;
  wire       [6:0]    _zz_refill_read_arbiter_oh_19;
  wire                _zz_refill_read_arbiter_oh_20;
  wire       [0:0]    _zz_refill_read_arbiter_oh_21;
  wire       [4:0]    _zz_refill_read_arbiter_oh_22;
  wire                _zz_refill_read_arbiter_oh_23;
  wire       [0:0]    _zz_refill_read_arbiter_oh_24;
  wire       [2:0]    _zz_refill_read_arbiter_oh_25;
  wire                _zz_refill_read_arbiter_oh_26;
  wire       [0:0]    _zz_refill_read_arbiter_oh_27;
  wire       [0:0]    _zz_refill_read_arbiter_oh_28;
  wire       [6:0]    _zz_refill_read_arbiter_oh_29;
  wire       [0:0]    _zz_refill_read_arbiter_oh_30;
  wire       [5:0]    _zz_refill_read_arbiter_oh_31;
  wire                _zz_refill_read_arbiter_oh_32;
  wire       [0:0]    _zz_refill_read_arbiter_oh_33;
  wire       [3:0]    _zz_refill_read_arbiter_oh_34;
  wire                _zz_refill_read_arbiter_oh_35;
  wire       [0:0]    _zz_refill_read_arbiter_oh_36;
  wire       [1:0]    _zz_refill_read_arbiter_oh_37;
  wire       [6:0]    _zz_refill_read_arbiter_oh_38;
  wire                _zz_refill_read_arbiter_oh_39;
  wire       [6:0]    _zz_refill_read_arbiter_oh_40;
  wire                _zz_refill_read_arbiter_oh_41;
  wire       [0:0]    _zz_refill_read_arbiter_oh_42;
  wire       [4:0]    _zz_refill_read_arbiter_oh_43;
  wire                _zz_refill_read_arbiter_oh_44;
  wire       [0:0]    _zz_refill_read_arbiter_oh_45;
  wire       [2:0]    _zz_refill_read_arbiter_oh_46;
  wire                _zz_refill_read_arbiter_oh_47;
  wire                _zz_refill_read_arbiter_oh_48;
  wire       [0:0]    _zz_refill_read_arbiter_oh_49;
  wire       [6:0]    _zz_refill_read_arbiter_oh_50;
  wire       [0:0]    _zz_refill_read_arbiter_oh_51;
  wire       [5:0]    _zz_refill_read_arbiter_oh_52;
  wire                _zz_refill_read_arbiter_oh_53;
  wire       [0:0]    _zz_refill_read_arbiter_oh_54;
  wire       [3:0]    _zz_refill_read_arbiter_oh_55;
  wire                _zz_refill_read_arbiter_oh_56;
  wire       [0:0]    _zz_refill_read_arbiter_oh_57;
  wire       [0:0]    _zz_refill_read_arbiter_oh_58;
  wire       [6:0]    _zz_refill_read_arbiter_oh_59;
  wire       [1:0]    _zz_refill_read_arbiter_oh_60;
  wire                _zz_refill_read_arbiter_oh_61;
  wire       [6:0]    _zz_refill_read_arbiter_oh_62;
  wire                _zz_refill_read_arbiter_oh_63;
  wire       [0:0]    _zz_refill_read_arbiter_oh_64;
  wire       [4:0]    _zz_refill_read_arbiter_oh_65;
  wire                _zz_refill_read_arbiter_oh_66;
  wire       [0:0]    _zz_refill_read_arbiter_oh_67;
  wire       [1:0]    _zz_refill_read_arbiter_oh_68;
  wire                _zz_refill_read_arbiter_oh_69;
  wire       [6:0]    _zz_refill_read_arbiter_oh_70;
  wire                _zz_refill_read_arbiter_oh_71;
  wire       [0:0]    _zz_refill_read_arbiter_oh_72;
  wire       [4:0]    _zz_refill_read_arbiter_oh_73;
  wire                _zz_refill_read_arbiter_oh_74;
  wire       [0:0]    _zz_refill_read_arbiter_oh_75;
  wire       [1:0]    _zz_refill_read_arbiter_oh_76;
  reg        [26:0]   _zz_refill_read_cmdAddress;
  reg        [31:0]   _zz_refill_read_rspAddress;
  reg        [0:0]    _zz_refill_read_way;
  wire       [7:0]    _zz__zz_writeback_free_1;
  wire                _zz_writeback_read_arbiter_oh;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_1;
  wire       [4:0]    _zz_writeback_read_arbiter_oh_2;
  wire                _zz_writeback_read_arbiter_oh_3;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_4;
  wire       [2:0]    _zz_writeback_read_arbiter_oh_5;
  wire                _zz_writeback_read_arbiter_oh_6;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_7;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_8;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_9;
  wire       [5:0]    _zz_writeback_read_arbiter_oh_10;
  wire                _zz_writeback_read_arbiter_oh_11;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_12;
  wire       [3:0]    _zz_writeback_read_arbiter_oh_13;
  wire                _zz_writeback_read_arbiter_oh_14;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_15;
  wire       [1:0]    _zz_writeback_read_arbiter_oh_16;
  wire                _zz_writeback_read_arbiter_oh_17;
  wire                _zz_writeback_read_arbiter_oh_18;
  wire       [6:0]    _zz_writeback_read_arbiter_oh_19;
  wire                _zz_writeback_read_arbiter_oh_20;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_21;
  wire       [4:0]    _zz_writeback_read_arbiter_oh_22;
  wire                _zz_writeback_read_arbiter_oh_23;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_24;
  wire       [2:0]    _zz_writeback_read_arbiter_oh_25;
  wire                _zz_writeback_read_arbiter_oh_26;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_27;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_28;
  wire       [6:0]    _zz_writeback_read_arbiter_oh_29;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_30;
  wire       [5:0]    _zz_writeback_read_arbiter_oh_31;
  wire                _zz_writeback_read_arbiter_oh_32;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_33;
  wire       [3:0]    _zz_writeback_read_arbiter_oh_34;
  wire                _zz_writeback_read_arbiter_oh_35;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_36;
  wire       [1:0]    _zz_writeback_read_arbiter_oh_37;
  wire       [6:0]    _zz_writeback_read_arbiter_oh_38;
  wire                _zz_writeback_read_arbiter_oh_39;
  wire       [6:0]    _zz_writeback_read_arbiter_oh_40;
  wire                _zz_writeback_read_arbiter_oh_41;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_42;
  wire       [4:0]    _zz_writeback_read_arbiter_oh_43;
  wire                _zz_writeback_read_arbiter_oh_44;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_45;
  wire       [2:0]    _zz_writeback_read_arbiter_oh_46;
  wire                _zz_writeback_read_arbiter_oh_47;
  wire                _zz_writeback_read_arbiter_oh_48;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_49;
  wire       [6:0]    _zz_writeback_read_arbiter_oh_50;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_51;
  wire       [5:0]    _zz_writeback_read_arbiter_oh_52;
  wire                _zz_writeback_read_arbiter_oh_53;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_54;
  wire       [3:0]    _zz_writeback_read_arbiter_oh_55;
  wire                _zz_writeback_read_arbiter_oh_56;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_57;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_58;
  wire       [6:0]    _zz_writeback_read_arbiter_oh_59;
  wire       [1:0]    _zz_writeback_read_arbiter_oh_60;
  wire                _zz_writeback_read_arbiter_oh_61;
  wire       [6:0]    _zz_writeback_read_arbiter_oh_62;
  wire                _zz_writeback_read_arbiter_oh_63;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_64;
  wire       [4:0]    _zz_writeback_read_arbiter_oh_65;
  wire                _zz_writeback_read_arbiter_oh_66;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_67;
  wire       [1:0]    _zz_writeback_read_arbiter_oh_68;
  wire                _zz_writeback_read_arbiter_oh_69;
  wire       [6:0]    _zz_writeback_read_arbiter_oh_70;
  wire                _zz_writeback_read_arbiter_oh_71;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_72;
  wire       [4:0]    _zz_writeback_read_arbiter_oh_73;
  wire                _zz_writeback_read_arbiter_oh_74;
  wire       [0:0]    _zz_writeback_read_arbiter_oh_75;
  wire       [1:0]    _zz_writeback_read_arbiter_oh_76;
  reg        [31:0]   _zz_writeback_read_address;
  reg        [0:0]    _zz_writeback_read_way;
  wire       [2:0]    _zz_writeback_read_wordIndex;
  wire       [0:0]    _zz_writeback_read_wordIndex_1;
  reg        [31:0]   _zz_writeback_read_readedData;
  wire       [5:0]    _zz_writeback_victimBuffer_port;
  wire                _zz_writeback_write_arbiter_oh;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_1;
  wire       [4:0]    _zz_writeback_write_arbiter_oh_2;
  wire                _zz_writeback_write_arbiter_oh_3;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_4;
  wire       [2:0]    _zz_writeback_write_arbiter_oh_5;
  wire                _zz_writeback_write_arbiter_oh_6;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_7;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_8;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_9;
  wire       [5:0]    _zz_writeback_write_arbiter_oh_10;
  wire                _zz_writeback_write_arbiter_oh_11;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_12;
  wire       [3:0]    _zz_writeback_write_arbiter_oh_13;
  wire                _zz_writeback_write_arbiter_oh_14;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_15;
  wire       [1:0]    _zz_writeback_write_arbiter_oh_16;
  wire                _zz_writeback_write_arbiter_oh_17;
  wire                _zz_writeback_write_arbiter_oh_18;
  wire       [6:0]    _zz_writeback_write_arbiter_oh_19;
  wire                _zz_writeback_write_arbiter_oh_20;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_21;
  wire       [4:0]    _zz_writeback_write_arbiter_oh_22;
  wire                _zz_writeback_write_arbiter_oh_23;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_24;
  wire       [2:0]    _zz_writeback_write_arbiter_oh_25;
  wire                _zz_writeback_write_arbiter_oh_26;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_27;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_28;
  wire       [6:0]    _zz_writeback_write_arbiter_oh_29;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_30;
  wire       [5:0]    _zz_writeback_write_arbiter_oh_31;
  wire                _zz_writeback_write_arbiter_oh_32;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_33;
  wire       [3:0]    _zz_writeback_write_arbiter_oh_34;
  wire                _zz_writeback_write_arbiter_oh_35;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_36;
  wire       [1:0]    _zz_writeback_write_arbiter_oh_37;
  wire       [6:0]    _zz_writeback_write_arbiter_oh_38;
  wire                _zz_writeback_write_arbiter_oh_39;
  wire       [6:0]    _zz_writeback_write_arbiter_oh_40;
  wire                _zz_writeback_write_arbiter_oh_41;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_42;
  wire       [4:0]    _zz_writeback_write_arbiter_oh_43;
  wire                _zz_writeback_write_arbiter_oh_44;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_45;
  wire       [2:0]    _zz_writeback_write_arbiter_oh_46;
  wire                _zz_writeback_write_arbiter_oh_47;
  wire                _zz_writeback_write_arbiter_oh_48;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_49;
  wire       [6:0]    _zz_writeback_write_arbiter_oh_50;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_51;
  wire       [5:0]    _zz_writeback_write_arbiter_oh_52;
  wire                _zz_writeback_write_arbiter_oh_53;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_54;
  wire       [3:0]    _zz_writeback_write_arbiter_oh_55;
  wire                _zz_writeback_write_arbiter_oh_56;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_57;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_58;
  wire       [6:0]    _zz_writeback_write_arbiter_oh_59;
  wire       [1:0]    _zz_writeback_write_arbiter_oh_60;
  wire                _zz_writeback_write_arbiter_oh_61;
  wire       [6:0]    _zz_writeback_write_arbiter_oh_62;
  wire                _zz_writeback_write_arbiter_oh_63;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_64;
  wire       [4:0]    _zz_writeback_write_arbiter_oh_65;
  wire                _zz_writeback_write_arbiter_oh_66;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_67;
  wire       [1:0]    _zz_writeback_write_arbiter_oh_68;
  wire                _zz_writeback_write_arbiter_oh_69;
  wire       [6:0]    _zz_writeback_write_arbiter_oh_70;
  wire                _zz_writeback_write_arbiter_oh_71;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_72;
  wire       [4:0]    _zz_writeback_write_arbiter_oh_73;
  wire                _zz_writeback_write_arbiter_oh_74;
  wire       [0:0]    _zz_writeback_write_arbiter_oh_75;
  wire       [1:0]    _zz_writeback_write_arbiter_oh_76;
  reg        [31:0]   _zz_writeback_write_bufferRead_payload_address;
  wire       [2:0]    _zz_writeback_write_wordIndex;
  wire       [0:0]    _zz_writeback_write_wordIndex_1;
  wire       [26:0]   _zz_load_pipeline_stages_1_REFILL_HITS_EARLY;
  wire       [26:0]   _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_1;
  wire                _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_2;
  wire                _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_3;
  wire       [0:0]    _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_4;
  wire       [1:0]    _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_5;
  reg                 _zz__zz_refill_push_payload_victim;
  reg                 _zz_load_ctrl_refillWayNeedWriteback;
  wire       [3:0]    _zz_load_ctrl_lineBusy;
  wire       [3:0]    _zz_load_ctrl_lineBusy_1;
  wire                _zz_load_ctrl_lineBusy_2;
  wire                _zz_load_ctrl_lineBusy_3;
  wire       [3:0]    _zz_load_ctrl_lineBusy_4;
  wire       [3:0]    _zz_load_ctrl_lineBusy_5;
  wire       [0:0]    _zz_load_ctrl_lineBusy_6;
  wire                _zz_load_ctrl_lineBusy_7;
  wire       [3:0]    _zz_load_ctrl_lineBusy_8;
  wire                _zz_load_ctrl_lineBusy_9;
  wire       [0:0]    _zz_load_ctrl_lineBusy_10;
  wire       [3:0]    _zz_load_ctrl_lineBusy_11;
  wire       [3:0]    _zz_load_ctrl_lineBusy_12;
  wire       [1:0]    _zz_load_ctrl_lineBusy_13;
  wire                _zz_load_ctrl_lineBusy_14;
  wire                _zz_load_ctrl_lineBusy_15;
  wire       [3:0]    _zz_load_ctrl_lineBusy_16;
  wire       [3:0]    _zz_load_ctrl_lineBusy_17;
  wire                _zz_load_ctrl_lineBusy_18;
  wire                _zz_load_ctrl_lineBusy_19;
  wire       [3:0]    _zz_load_ctrl_lineBusy_20;
  wire       [3:0]    _zz_load_ctrl_lineBusy_21;
  wire       [0:0]    _zz_load_ctrl_lineBusy_22;
  wire                _zz_load_ctrl_lineBusy_23;
  wire       [3:0]    _zz_load_ctrl_lineBusy_24;
  wire                _zz_load_ctrl_lineBusy_25;
  wire       [0:0]    _zz_load_ctrl_lineBusy_26;
  wire       [3:0]    _zz_load_ctrl_lineBusy_27;
  wire       [3:0]    _zz_load_ctrl_lineBusy_28;
  wire       [1:0]    _zz_load_ctrl_lineBusy_29;
  wire                _zz_load_ctrl_lineBusy_30;
  wire                _zz_load_ctrl_lineBusy_31;
  reg        [22:0]   _zz_writeback_push_payload_address;
  wire       [26:0]   _zz_store_pipeline_stages_1_REFILL_HITS_EARLY;
  wire       [26:0]   _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_1;
  wire                _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_2;
  wire                _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_3;
  wire       [0:0]    _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_4;
  wire       [1:0]    _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_5;
  reg                 _zz_store_ctrl_replacedWayNeedWriteback;
  reg                 _zz_store_ctrl_replacedWayNeedWriteback_1;
  wire       [3:0]    _zz_store_ctrl_lineBusy;
  wire       [3:0]    _zz_store_ctrl_lineBusy_1;
  wire                _zz_store_ctrl_lineBusy_2;
  wire                _zz_store_ctrl_lineBusy_3;
  wire       [3:0]    _zz_store_ctrl_lineBusy_4;
  wire       [3:0]    _zz_store_ctrl_lineBusy_5;
  wire       [0:0]    _zz_store_ctrl_lineBusy_6;
  wire                _zz_store_ctrl_lineBusy_7;
  wire       [3:0]    _zz_store_ctrl_lineBusy_8;
  wire                _zz_store_ctrl_lineBusy_9;
  wire       [0:0]    _zz_store_ctrl_lineBusy_10;
  wire       [3:0]    _zz_store_ctrl_lineBusy_11;
  wire       [3:0]    _zz_store_ctrl_lineBusy_12;
  wire       [1:0]    _zz_store_ctrl_lineBusy_13;
  wire                _zz_store_ctrl_lineBusy_14;
  wire                _zz_store_ctrl_lineBusy_15;
  wire       [3:0]    _zz_store_ctrl_lineBusy_16;
  wire       [3:0]    _zz_store_ctrl_lineBusy_17;
  wire                _zz_store_ctrl_lineBusy_18;
  wire                _zz_store_ctrl_lineBusy_19;
  wire       [3:0]    _zz_store_ctrl_lineBusy_20;
  wire       [3:0]    _zz_store_ctrl_lineBusy_21;
  wire       [0:0]    _zz_store_ctrl_lineBusy_22;
  wire                _zz_store_ctrl_lineBusy_23;
  wire       [3:0]    _zz_store_ctrl_lineBusy_24;
  wire                _zz_store_ctrl_lineBusy_25;
  wire       [0:0]    _zz_store_ctrl_lineBusy_26;
  wire       [3:0]    _zz_store_ctrl_lineBusy_27;
  wire       [3:0]    _zz_store_ctrl_lineBusy_28;
  wire       [1:0]    _zz_store_ctrl_lineBusy_29;
  wire                _zz_store_ctrl_lineBusy_30;
  wire                _zz_store_ctrl_lineBusy_31;
  reg        [22:0]   _zz_writeback_push_payload_address_1;
  reg                 _zz_refill_push_payload_victim_1;
  wire       [0:0]    _zz_when;
  wire       [0:0]    _zz_when_1;
  wire                store_pipeline_stages_0_isThrown;
  wire                store_pipeline_stages_1_isThrown;
  wire                store_pipeline_stages_2_isThrown;
  reg        [2:0]    store_pipeline_stages_1_TRANSACTION_ID;
  reg                 store_pipeline_stages_1_FLUSH_FREE;
  reg        [3:0]    store_pipeline_stages_1_CPU_MASK;
  reg        [31:0]   store_pipeline_stages_1_CPU_WORD;
  reg                 store_pipeline_stages_1_IO;
  reg                 store_pipeline_stages_1_PREFETCH;
  reg                 store_pipeline_stages_1_FLUSH;
  reg        [2:0]    store_pipeline_stages_2_TRANSACTION_ID;
  reg                 store_pipeline_stages_2_FLUSH_FREE;
  reg        [3:0]    store_pipeline_stages_2_CPU_MASK;
  reg        [31:0]   store_pipeline_stages_2_CPU_WORD;
  reg                 store_pipeline_stages_2_IO;
  wire       [7:0]    store_pipeline_stages_2_REFILL_SLOT;
  wire                store_pipeline_stages_2_REFILL_SLOT_FULL;
  reg                 store_pipeline_stages_2_WAYS_HIT;
  reg                 store_pipeline_stages_2_MISS;
  reg                 store_pipeline_stages_2_REDO;
  reg                 store_pipeline_stages_2_PREFETCH;
  reg                 store_pipeline_stages_2_FLUSH;
  wire       [1:0]    store_pipeline_stages_2_WAYS_HAZARD_resulting;
  reg        [1:0]    store_pipeline_stages_2_WAYS_HITS;
  reg                 store_pipeline_stages_2_STATUS_0_dirty;
  reg                 store_pipeline_stages_2_STATUS_1_dirty;
  reg                 store_pipeline_stages_2_WAYS_TAGS_0_loaded;
  reg        [22:0]   store_pipeline_stages_2_WAYS_TAGS_0_address;
  reg                 store_pipeline_stages_2_WAYS_TAGS_0_fault;
  reg                 store_pipeline_stages_2_WAYS_TAGS_1_loaded;
  reg        [22:0]   store_pipeline_stages_2_WAYS_TAGS_1_address;
  reg                 store_pipeline_stages_2_WAYS_TAGS_1_fault;
  reg        [7:0]    store_pipeline_stages_2_REFILL_HITS_EARLY;
  wire       [7:0]    store_pipeline_stages_2_REFILL_HITS;
  reg        [7:0]    store_pipeline_stages_1_REFILL_HITS_EARLY;
  wire                store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  wire                store_pipeline_stages_1_STATUS_overloaded_1_dirty;
  wire                store_pipeline_stages_1_STATUS_0_dirty;
  wire                store_pipeline_stages_1_STATUS_1_dirty;
  wire                store_pipeline_stages_1_WAYS_HIT;
  reg        [1:0]    store_pipeline_stages_1_WAYS_HITS;
  wire                store_pipeline_stages_1_WAYS_TAGS_0_loaded;
  wire       [22:0]   store_pipeline_stages_1_WAYS_TAGS_0_address;
  wire                store_pipeline_stages_1_WAYS_TAGS_0_fault;
  wire                store_pipeline_stages_1_WAYS_TAGS_1_loaded;
  wire       [22:0]   store_pipeline_stages_1_WAYS_TAGS_1_address;
  wire                store_pipeline_stages_1_WAYS_TAGS_1_fault;
  wire                store_pipeline_stages_1_ready;
  wire       [1:0]    store_pipeline_stages_0_WAYS_HAZARD;
  wire       [2:0]    store_pipeline_stages_0_TRANSACTION_ID;
  wire                store_pipeline_stages_0_PREFETCH;
  wire                store_pipeline_stages_0_FLUSH_FREE;
  wire                store_pipeline_stages_0_FLUSH;
  wire                store_pipeline_stages_0_IO;
  wire       [3:0]    store_pipeline_stages_0_CPU_MASK;
  wire       [31:0]   store_pipeline_stages_0_CPU_WORD;
  wire       [31:0]   store_pipeline_stages_0_ADDRESS_POST_TRANSLATION;
  reg        [31:0]   store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  reg        [1:0]    store_pipeline_stages_2_WAYS_HAZARD;
  wire       [1:0]    store_pipeline_stages_2_WAYS_HAZARD_overloaded;
  reg        [31:0]   store_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
  reg        [1:0]    store_pipeline_stages_1_WAYS_HAZARD;
  wire       [1:0]    store_pipeline_stages_1_WAYS_HAZARD_overloaded;
  wire                load_pipeline_stages_0_isThrown;
  wire                load_pipeline_stages_1_isThrown;
  wire                load_pipeline_stages_2_isThrown;
  reg        [2:0]    load_pipeline_stages_1_TRANSACTION_ID;
  reg                 load_pipeline_stages_1_ABORD;
  reg        [1:0]    load_pipeline_stages_2_WAYS_HAZARD;
  reg        [2:0]    load_pipeline_stages_2_TRANSACTION_ID;
  wire       [7:0]    load_pipeline_stages_2_REFILL_SLOT;
  wire                load_pipeline_stages_2_REFILL_SLOT_FULL;
  reg                 load_pipeline_stages_2_ABORD;
  wire                load_pipeline_stages_2_FAULT;
  reg                 load_pipeline_stages_2_MISS;
  reg                 load_pipeline_stages_2_REDO;
  wire       [1:0]    load_pipeline_stages_2_WAYS_HAZARD_resulting;
  reg        [1:0]    load_pipeline_stages_2_BANK_BUSY_REMAPPED;
  reg        [31:0]   load_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  reg                 load_pipeline_stages_2_STATUS_0_dirty;
  reg                 load_pipeline_stages_2_STATUS_1_dirty;
  reg                 load_pipeline_stages_2_WAYS_TAGS_0_loaded;
  reg        [22:0]   load_pipeline_stages_2_WAYS_TAGS_0_address;
  reg                 load_pipeline_stages_2_WAYS_TAGS_0_fault;
  reg                 load_pipeline_stages_2_WAYS_TAGS_1_loaded;
  reg        [22:0]   load_pipeline_stages_2_WAYS_TAGS_1_address;
  reg                 load_pipeline_stages_2_WAYS_TAGS_1_fault;
  reg        [7:0]    load_pipeline_stages_2_REFILL_HITS_EARLY;
  wire       [7:0]    load_pipeline_stages_2_REFILL_HITS;
  reg        [7:0]    load_pipeline_stages_1_REFILL_HITS_EARLY;
  wire                load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  wire                load_pipeline_stages_1_STATUS_overloaded_1_dirty;
  wire                load_pipeline_stages_1_STATUS_0_dirty;
  wire                load_pipeline_stages_1_STATUS_1_dirty;
  wire                load_pipeline_stages_2_WAYS_HIT;
  reg        [31:0]   load_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
  reg        [1:0]    load_pipeline_stages_1_WAYS_HITS;
  wire                load_pipeline_stages_1_WAYS_TAGS_0_loaded;
  wire       [22:0]   load_pipeline_stages_1_WAYS_TAGS_0_address;
  wire                load_pipeline_stages_1_WAYS_TAGS_0_fault;
  wire                load_pipeline_stages_1_WAYS_TAGS_1_loaded;
  wire       [22:0]   load_pipeline_stages_1_WAYS_TAGS_1_address;
  wire                load_pipeline_stages_1_WAYS_TAGS_1_fault;
  wire                load_pipeline_stages_1_ready;
  wire                load_pipeline_stages_0_ABORD;
  wire       [31:0]   load_pipeline_stages_0_ADDRESS_POST_TRANSLATION;
  reg        [31:0]   load_pipeline_stages_2_BANKS_MUXES_0;
  reg        [31:0]   load_pipeline_stages_2_BANKS_MUXES_1;
  reg        [1:0]    load_pipeline_stages_2_WAYS_HITS;
  wire       [31:0]   load_pipeline_stages_2_CPU_WORD;
  wire       [31:0]   load_pipeline_stages_1_BANKS_MUXES_0;
  wire       [31:0]   load_pipeline_stages_1_BANKS_MUXES_1;
  reg        [1:0]    load_pipeline_stages_1_BANK_BUSY;
  reg        [1:0]    load_pipeline_stages_1_BANK_BUSY_REMAPPED;
  wire       [31:0]   load_pipeline_stages_1_BANKS_WORDS_0;
  wire       [31:0]   load_pipeline_stages_1_BANKS_WORDS_1;
  reg        [1:0]    load_pipeline_stages_0_BANK_BUSY_overloaded;
  wire                load_pipeline_stages_0_ready;
  reg        [1:0]    load_pipeline_stages_0_BANK_BUSY;
  wire       [1:0]    load_pipeline_stages_0_WAYS_HAZARD;
  wire       [2:0]    load_pipeline_stages_0_TRANSACTION_ID;
  wire                load_pipeline_stages_0_REDO_ON_DATA_HAZARD;
  wire       [31:0]   load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION;
  reg        [31:0]   load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION;
  reg        [1:0]    load_pipeline_stages_1_WAYS_HAZARD;
  wire       [1:0]    load_pipeline_stages_1_WAYS_HAZARD_overloaded;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 banks_0_write_valid;
  reg        [6:0]    banks_0_write_payload_address;
  reg        [31:0]   banks_0_write_payload_data;
  reg        [3:0]    banks_0_write_payload_mask;
  reg                 banks_0_read_usedByWriteBack;
  reg                 banks_0_read_cmd_valid;
  reg        [6:0]    banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [31:0]   banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  reg                 banks_1_write_valid;
  reg        [6:0]    banks_1_write_payload_address;
  reg        [31:0]   banks_1_write_payload_data;
  reg        [3:0]    banks_1_write_payload_mask;
  reg                 banks_1_read_usedByWriteBack;
  reg                 banks_1_read_cmd_valid;
  reg        [6:0]    banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [31:0]   banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [1:0]    waysWrite_mask;
  reg        [3:0]    waysWrite_address;
  reg                 waysWrite_tag_loaded;
  reg        [22:0]   waysWrite_tag_address;
  reg                 waysWrite_tag_fault;
  reg        [1:0]    waysWrite_maskLast;
  reg        [3:0]    waysWrite_addressLast;
  wire                ways_0_loadRead_cmd_valid;
  wire       [3:0]    ways_0_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_0_loadRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [22:0]   ways_0_loadRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_0_loadRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [24:0]   _zz_ways_0_loadRead_rsp_loaded;
  wire                ways_0_storeRead_cmd_valid;
  wire       [3:0]    ways_0_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_0_storeRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [22:0]   ways_0_storeRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_0_storeRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [24:0]   _zz_ways_0_storeRead_rsp_loaded;
  wire                ways_1_loadRead_cmd_valid;
  wire       [3:0]    ways_1_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_1_loadRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [22:0]   ways_1_loadRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_1_loadRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [24:0]   _zz_ways_1_loadRead_rsp_loaded;
  wire                ways_1_storeRead_cmd_valid;
  wire       [3:0]    ways_1_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_1_storeRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [22:0]   ways_1_storeRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_1_storeRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [24:0]   _zz_ways_1_storeRead_rsp_loaded;
  reg                 status_write_valid;
  reg        [3:0]    status_write_payload_address;
  reg                 status_write_payload_data_0_dirty;
  reg                 status_write_payload_data_1_dirty;
  wire                status_loadRead_cmd_valid;
  wire       [3:0]    status_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                status_loadRead_rsp_0_dirty /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                status_loadRead_rsp_1_dirty /* synthesis syn_keep = 1 */ ;
  wire       [1:0]    _zz_status_loadRead_rsp_0_dirty;
  wire                status_storeRead_cmd_valid;
  wire       [3:0]    status_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                status_storeRead_rsp_0_dirty /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                status_storeRead_rsp_1_dirty /* synthesis syn_keep = 1 */ ;
  wire       [1:0]    _zz_status_storeRead_rsp_0_dirty;
  reg                 status_writeLast_valid;
  reg        [3:0]    status_writeLast_payload_address;
  reg                 status_writeLast_payload_data_0_dirty;
  reg                 status_writeLast_payload_data_1_dirty;
  wire                wayRandom_willIncrement;
  wire                wayRandom_willClear;
  reg        [0:0]    wayRandom_valueNext;
  reg        [0:0]    wayRandom_value;
  wire                wayRandom_willOverflowIfInc;
  wire                wayRandom_willOverflow;
  reg        [4:0]    invalidate_counter;
  wire                invalidate_done;
  wire                invalidate_reservation_win;
  reg                 invalidate_reservation_take;
  wire                when_dcache2_l680;
  reg                 invalidate_done_regNext;
  reg                 refill_slots_0_valid;
  reg        [31:0]   refill_slots_0_address;
  reg        [0:0]    refill_slots_0_way;
  reg                 refill_slots_0_cmdSent;
  reg        [6:0]    refill_slots_0_priority;
  reg                 refill_slots_0_loaded;
  reg        [0:0]    refill_slots_0_loadedCounter;
  wire                refill_slots_0_loadedDone;
  wire                refill_slots_0_free;
  reg        [7:0]    refill_slots_0_victim;
  reg        [7:0]    refill_slots_0_writebackHazards;
  reg                 refill_slots_1_valid;
  reg        [31:0]   refill_slots_1_address;
  reg        [0:0]    refill_slots_1_way;
  reg                 refill_slots_1_cmdSent;
  reg        [6:0]    refill_slots_1_priority;
  reg                 refill_slots_1_loaded;
  reg        [0:0]    refill_slots_1_loadedCounter;
  wire                refill_slots_1_loadedDone;
  wire                refill_slots_1_free;
  reg        [7:0]    refill_slots_1_victim;
  reg        [7:0]    refill_slots_1_writebackHazards;
  reg                 refill_slots_2_valid;
  reg        [31:0]   refill_slots_2_address;
  reg        [0:0]    refill_slots_2_way;
  reg                 refill_slots_2_cmdSent;
  reg        [6:0]    refill_slots_2_priority;
  reg                 refill_slots_2_loaded;
  reg        [0:0]    refill_slots_2_loadedCounter;
  wire                refill_slots_2_loadedDone;
  wire                refill_slots_2_free;
  reg        [7:0]    refill_slots_2_victim;
  reg        [7:0]    refill_slots_2_writebackHazards;
  reg                 refill_slots_3_valid;
  reg        [31:0]   refill_slots_3_address;
  reg        [0:0]    refill_slots_3_way;
  reg                 refill_slots_3_cmdSent;
  reg        [6:0]    refill_slots_3_priority;
  reg                 refill_slots_3_loaded;
  reg        [0:0]    refill_slots_3_loadedCounter;
  wire                refill_slots_3_loadedDone;
  wire                refill_slots_3_free;
  reg        [7:0]    refill_slots_3_victim;
  reg        [7:0]    refill_slots_3_writebackHazards;
  reg                 refill_slots_4_valid;
  reg        [31:0]   refill_slots_4_address;
  reg        [0:0]    refill_slots_4_way;
  reg                 refill_slots_4_cmdSent;
  reg        [6:0]    refill_slots_4_priority;
  reg                 refill_slots_4_loaded;
  reg        [0:0]    refill_slots_4_loadedCounter;
  wire                refill_slots_4_loadedDone;
  wire                refill_slots_4_free;
  reg        [7:0]    refill_slots_4_victim;
  reg        [7:0]    refill_slots_4_writebackHazards;
  reg                 refill_slots_5_valid;
  reg        [31:0]   refill_slots_5_address;
  reg        [0:0]    refill_slots_5_way;
  reg                 refill_slots_5_cmdSent;
  reg        [6:0]    refill_slots_5_priority;
  reg                 refill_slots_5_loaded;
  reg        [0:0]    refill_slots_5_loadedCounter;
  wire                refill_slots_5_loadedDone;
  wire                refill_slots_5_free;
  reg        [7:0]    refill_slots_5_victim;
  reg        [7:0]    refill_slots_5_writebackHazards;
  reg                 refill_slots_6_valid;
  reg        [31:0]   refill_slots_6_address;
  reg        [0:0]    refill_slots_6_way;
  reg                 refill_slots_6_cmdSent;
  reg        [6:0]    refill_slots_6_priority;
  reg                 refill_slots_6_loaded;
  reg        [0:0]    refill_slots_6_loadedCounter;
  wire                refill_slots_6_loadedDone;
  wire                refill_slots_6_free;
  reg        [7:0]    refill_slots_6_victim;
  reg        [7:0]    refill_slots_6_writebackHazards;
  reg                 refill_slots_7_valid;
  reg        [31:0]   refill_slots_7_address;
  reg        [0:0]    refill_slots_7_way;
  reg                 refill_slots_7_cmdSent;
  reg        [6:0]    refill_slots_7_priority;
  reg                 refill_slots_7_loaded;
  reg        [0:0]    refill_slots_7_loadedCounter;
  wire                refill_slots_7_loadedDone;
  wire                refill_slots_7_free;
  reg        [7:0]    refill_slots_7_victim;
  reg        [7:0]    refill_slots_7_writebackHazards;
  wire       [7:0]    _zz_refill_free;
  wire       [7:0]    _zz_refill_free_1;
  wire       [7:0]    refill_free;
  wire                refill_full;
  reg                 refill_push_valid;
  reg        [31:0]   refill_push_payload_address;
  reg        [0:0]    refill_push_payload_way;
  reg        [7:0]    refill_push_payload_victim;
  wire                when_dcache2_l750;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                when_dcache2_l750_1;
  wire                when_dcache2_l750_2;
  wire                when_dcache2_l750_3;
  wire                when_dcache2_l750_4;
  wire                when_dcache2_l750_5;
  wire                when_dcache2_l750_6;
  wire                when_dcache2_l750_7;
  wire                refill_read_arbiter_slotsWithId_0_0;
  wire                refill_read_arbiter_slotsWithId_1_0;
  wire                refill_read_arbiter_slotsWithId_2_0;
  wire                refill_read_arbiter_slotsWithId_3_0;
  wire                refill_read_arbiter_slotsWithId_4_0;
  wire                refill_read_arbiter_slotsWithId_5_0;
  wire                refill_read_arbiter_slotsWithId_6_0;
  wire                refill_read_arbiter_slotsWithId_7_0;
  wire       [7:0]    refill_read_arbiter_hits;
  wire                refill_read_arbiter_hit;
  reg        [7:0]    refill_read_arbiter_oh;
  wire                _zz_refill_read_arbiter_sel;
  wire                _zz_refill_read_arbiter_sel_1;
  wire                _zz_refill_read_arbiter_sel_2;
  wire                _zz_refill_read_arbiter_sel_3;
  wire                _zz_refill_read_arbiter_sel_4;
  wire                _zz_refill_read_arbiter_sel_5;
  wire                _zz_refill_read_arbiter_sel_6;
  wire                _zz_refill_read_arbiter_sel_7;
  wire                _zz_refill_read_arbiter_sel_8;
  wire                _zz_refill_read_arbiter_sel_9;
  wire       [2:0]    refill_read_arbiter_sel;
  reg        [7:0]    refill_read_arbiter_lock;
  wire                when_dcache2_l707;
  reg        [7:0]    refill_read_writebackHazards;
  wire                refill_read_writebackHazard;
  wire                io_mem_read_cmd_fire;
  wire                when_dcache2_l779;
  wire       [31:0]   refill_read_cmdAddress;
  wire                when_dcache2_l791;
  wire                when_dcache2_l791_1;
  wire                when_dcache2_l791_2;
  wire                when_dcache2_l791_3;
  wire                when_dcache2_l791_4;
  wire                when_dcache2_l791_5;
  wire                when_dcache2_l791_6;
  wire                when_dcache2_l791_7;
  wire       [31:0]   refill_read_rspAddress;
  wire       [0:0]    refill_read_way;
  (* keep , syn_keep *) reg        [2:0]    refill_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                refill_read_rspWithData;
  reg        [1:0]    refill_read_bankWriteNotif;
  reg                 refill_read_hadError;
  wire                when_dcache2_l821;
  reg                 refill_read_fire;
  wire                refill_read_reservation_win;
  reg                 refill_read_reservation_take;
  wire                refill_read_faulty;
  wire                when_dcache2_l834;
  reg                 writeback_slots_0_fire;
  reg                 writeback_slots_0_valid;
  reg        [31:0]   writeback_slots_0_address;
  reg        [0:0]    writeback_slots_0_way;
  reg        [6:0]    writeback_slots_0_priority;
  reg                 writeback_slots_0_readCmdDone;
  reg                 writeback_slots_0_victimBufferReady;
  reg                 writeback_slots_0_readRspDone;
  reg                 writeback_slots_0_writeCmdDone;
  wire                writeback_slots_0_free;
  reg                 writeback_slots_1_fire;
  reg                 writeback_slots_1_valid;
  reg        [31:0]   writeback_slots_1_address;
  reg        [0:0]    writeback_slots_1_way;
  reg        [6:0]    writeback_slots_1_priority;
  reg                 writeback_slots_1_readCmdDone;
  reg                 writeback_slots_1_victimBufferReady;
  reg                 writeback_slots_1_readRspDone;
  reg                 writeback_slots_1_writeCmdDone;
  wire                writeback_slots_1_free;
  reg                 writeback_slots_2_fire;
  reg                 writeback_slots_2_valid;
  reg        [31:0]   writeback_slots_2_address;
  reg        [0:0]    writeback_slots_2_way;
  reg        [6:0]    writeback_slots_2_priority;
  reg                 writeback_slots_2_readCmdDone;
  reg                 writeback_slots_2_victimBufferReady;
  reg                 writeback_slots_2_readRspDone;
  reg                 writeback_slots_2_writeCmdDone;
  wire                writeback_slots_2_free;
  reg                 writeback_slots_3_fire;
  reg                 writeback_slots_3_valid;
  reg        [31:0]   writeback_slots_3_address;
  reg        [0:0]    writeback_slots_3_way;
  reg        [6:0]    writeback_slots_3_priority;
  reg                 writeback_slots_3_readCmdDone;
  reg                 writeback_slots_3_victimBufferReady;
  reg                 writeback_slots_3_readRspDone;
  reg                 writeback_slots_3_writeCmdDone;
  wire                writeback_slots_3_free;
  reg                 writeback_slots_4_fire;
  reg                 writeback_slots_4_valid;
  reg        [31:0]   writeback_slots_4_address;
  reg        [0:0]    writeback_slots_4_way;
  reg        [6:0]    writeback_slots_4_priority;
  reg                 writeback_slots_4_readCmdDone;
  reg                 writeback_slots_4_victimBufferReady;
  reg                 writeback_slots_4_readRspDone;
  reg                 writeback_slots_4_writeCmdDone;
  wire                writeback_slots_4_free;
  reg                 writeback_slots_5_fire;
  reg                 writeback_slots_5_valid;
  reg        [31:0]   writeback_slots_5_address;
  reg        [0:0]    writeback_slots_5_way;
  reg        [6:0]    writeback_slots_5_priority;
  reg                 writeback_slots_5_readCmdDone;
  reg                 writeback_slots_5_victimBufferReady;
  reg                 writeback_slots_5_readRspDone;
  reg                 writeback_slots_5_writeCmdDone;
  wire                writeback_slots_5_free;
  reg                 writeback_slots_6_fire;
  reg                 writeback_slots_6_valid;
  reg        [31:0]   writeback_slots_6_address;
  reg        [0:0]    writeback_slots_6_way;
  reg        [6:0]    writeback_slots_6_priority;
  reg                 writeback_slots_6_readCmdDone;
  reg                 writeback_slots_6_victimBufferReady;
  reg                 writeback_slots_6_readRspDone;
  reg                 writeback_slots_6_writeCmdDone;
  wire                writeback_slots_6_free;
  reg                 writeback_slots_7_fire;
  reg                 writeback_slots_7_valid;
  reg        [31:0]   writeback_slots_7_address;
  reg        [0:0]    writeback_slots_7_way;
  reg        [6:0]    writeback_slots_7_priority;
  reg                 writeback_slots_7_readCmdDone;
  reg                 writeback_slots_7_victimBufferReady;
  reg                 writeback_slots_7_readRspDone;
  reg                 writeback_slots_7_writeCmdDone;
  wire                writeback_slots_7_free;
  wire       [7:0]    _zz_writeback_free;
  wire       [7:0]    _zz_writeback_free_1;
  wire       [7:0]    writeback_free;
  wire                writeback_full;
  reg                 writeback_push_valid;
  reg        [31:0]   writeback_push_payload_address;
  reg        [0:0]    writeback_push_payload_way;
  wire                when_dcache2_l897;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                when_dcache2_l897_1;
  wire                when_dcache2_l897_2;
  wire                when_dcache2_l897_3;
  wire                when_dcache2_l897_4;
  wire                when_dcache2_l897_5;
  wire                when_dcache2_l897_6;
  wire                when_dcache2_l897_7;
  wire                writeback_read_arbiter_slotsWithId_0_0;
  wire                writeback_read_arbiter_slotsWithId_1_0;
  wire                writeback_read_arbiter_slotsWithId_2_0;
  wire                writeback_read_arbiter_slotsWithId_3_0;
  wire                writeback_read_arbiter_slotsWithId_4_0;
  wire                writeback_read_arbiter_slotsWithId_5_0;
  wire                writeback_read_arbiter_slotsWithId_6_0;
  wire                writeback_read_arbiter_slotsWithId_7_0;
  wire       [7:0]    writeback_read_arbiter_hits;
  wire                writeback_read_arbiter_hit;
  reg        [7:0]    writeback_read_arbiter_oh;
  wire                _zz_writeback_read_arbiter_sel;
  wire                _zz_writeback_read_arbiter_sel_1;
  wire                _zz_writeback_read_arbiter_sel_2;
  wire                _zz_writeback_read_arbiter_sel_3;
  wire                _zz_writeback_read_arbiter_sel_4;
  wire                _zz_writeback_read_arbiter_sel_5;
  wire                _zz_writeback_read_arbiter_sel_6;
  wire                _zz_writeback_read_arbiter_sel_7;
  wire                _zz_writeback_read_arbiter_sel_8;
  wire                _zz_writeback_read_arbiter_sel_9;
  wire       [2:0]    writeback_read_arbiter_sel;
  reg        [7:0]    writeback_read_arbiter_lock;
  wire                when_dcache2_l707_1;
  wire       [31:0]   writeback_read_address;
  wire       [0:0]    writeback_read_way;
  (* keep , syn_keep *) reg        [2:0]    writeback_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                writeback_read_slotRead_valid;
  wire       [2:0]    writeback_read_slotRead_payload_id;
  wire                writeback_read_slotRead_payload_last;
  wire       [2:0]    writeback_read_slotRead_payload_wordIndex;
  wire       [0:0]    writeback_read_slotRead_payload_way;
  wire                when_dcache2_l937;
  wire                when_dcache2_l948;
  wire                when_dcache2_l948_1;
  reg                 writeback_read_slotReadLast_valid;
  reg        [2:0]    writeback_read_slotReadLast_payload_id;
  reg                 writeback_read_slotReadLast_payload_last;
  reg        [2:0]    writeback_read_slotReadLast_payload_wordIndex;
  reg        [0:0]    writeback_read_slotReadLast_payload_way;
  wire       [31:0]   writeback_read_readedData;
  wire                writeback_write_arbiter_slotsWithId_0_0;
  wire                writeback_write_arbiter_slotsWithId_1_0;
  wire                writeback_write_arbiter_slotsWithId_2_0;
  wire                writeback_write_arbiter_slotsWithId_3_0;
  wire                writeback_write_arbiter_slotsWithId_4_0;
  wire                writeback_write_arbiter_slotsWithId_5_0;
  wire                writeback_write_arbiter_slotsWithId_6_0;
  wire                writeback_write_arbiter_slotsWithId_7_0;
  wire       [7:0]    writeback_write_arbiter_hits;
  wire                writeback_write_arbiter_hit;
  reg        [7:0]    writeback_write_arbiter_oh;
  wire                _zz_writeback_write_arbiter_sel;
  wire                _zz_writeback_write_arbiter_sel_1;
  wire                _zz_writeback_write_arbiter_sel_2;
  wire                _zz_writeback_write_arbiter_sel_3;
  wire                _zz_writeback_write_arbiter_sel_4;
  wire                _zz_writeback_write_arbiter_sel_5;
  wire                _zz_writeback_write_arbiter_sel_6;
  wire                _zz_writeback_write_arbiter_sel_7;
  wire                _zz_writeback_write_arbiter_sel_8;
  wire                _zz_writeback_write_arbiter_sel_9;
  wire       [2:0]    writeback_write_arbiter_sel;
  reg        [7:0]    writeback_write_arbiter_lock;
  wire                when_dcache2_l707_2;
  (* keep , syn_keep *) reg        [2:0]    writeback_write_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                writeback_write_last;
  wire                writeback_write_bufferRead_valid;
  reg                 writeback_write_bufferRead_ready;
  wire       [2:0]    writeback_write_bufferRead_payload_id;
  wire       [31:0]   writeback_write_bufferRead_payload_address;
  wire                writeback_write_bufferRead_payload_last;
  wire                writeback_write_bufferRead_fire;
  wire                when_dcache2_l1020;
  wire                writeback_write_cmd_valid;
  wire                writeback_write_cmd_ready;
  wire       [2:0]    writeback_write_cmd_payload_id;
  wire       [31:0]   writeback_write_cmd_payload_address;
  wire                writeback_write_cmd_payload_last;
  reg                 writeback_write_bufferRead_rValid;
  reg        [2:0]    writeback_write_bufferRead_rData_id;
  reg        [31:0]   writeback_write_bufferRead_rData_address;
  reg                 writeback_write_bufferRead_rData_last;
  wire                when_Stream_l477;
  wire       [5:0]    _zz_writeback_write_word;
  wire       [31:0]   writeback_write_word;
  wire                load_pipeline_stages_0_valid;
  reg                 _zz_load_pipeline_stages_1_valid;
  reg                 load_pipeline_stages_1_valid;
  reg                 _zz_load_pipeline_stages_2_valid;
  reg                 load_pipeline_stages_2_valid;
  wire                _zz_load_pipeline_stages_0_throwRequest_dcache2_l1064;
  wire                load_pipeline_stages_0_throwRequest_dcache2_l1064;
  wire                _zz_load_pipeline_stages_1_throwRequest_dcache2_l1064;
  wire                load_pipeline_stages_1_throwRequest_dcache2_l1064;
  wire                load_pipeline_stages_2_throwRequest_dcache2_l1064;
  wire                when_dcache2_l1108;
  wire                when_dcache2_l1108_1;
  wire                _zz_load_pipeline_stages_2_CPU_WORD;
  reg                 _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  reg                 _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty;
  wire                when_dcache2_l659;
  wire                when_dcache2_l662;
  wire                load_refillCheckEarly_refillPushHit;
  wire                load_ctrl_reservation_win;
  reg                 load_ctrl_reservation_take;
  wire       [0:0]    load_ctrl_refillWay;
  wire                _zz_refill_push_payload_victim;
  wire                load_ctrl_refillWayNeedWriteback;
  wire                load_ctrl_refillHit;
  wire                load_ctrl_refillLoaded;
  wire                load_ctrl_lineBusy;
  wire                load_ctrl_bankBusy;
  wire                load_ctrl_waysHitHazard;
  wire                load_ctrl_canRefill;
  wire                load_ctrl_askRefill;
  wire                load_ctrl_startRefill;
  wire       [0:0]    load_ctrl_wayId;
  wire       [1:0]    _zz_34;
  wire                when_Pipeline_l276;
  wire                when_Pipeline_l276_1;
  wire                store_pipeline_stages_0_valid;
  reg                 _zz_store_pipeline_stages_1_valid;
  reg                 store_pipeline_stages_1_valid;
  reg                 _zz_store_pipeline_stages_2_valid;
  reg                 store_pipeline_stages_2_valid;
  wire                store_pipeline_discardAll;
  wire                store_pipeline_stages_0_throwRequest_dcache2_l1357;
  wire                store_pipeline_stages_1_throwRequest_dcache2_l1357;
  wire                store_pipeline_stages_2_throwRequest_dcache2_l1357;
  wire                _zz_35;
  wire                _zz_36;
  wire       [0:0]    _zz_37;
  wire       [1:0]    _zz_38;
  reg                 _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  reg                 _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty;
  wire                when_dcache2_l659_1;
  wire                when_dcache2_l662_1;
  wire                store_refillCheckEarly_refillPushHit;
  wire                store_ctrl_generationOk;
  wire                store_ctrl_reservation_win;
  reg                 store_ctrl_reservation_take;
  wire       [0:0]    store_ctrl_replacedWay;
  wire                store_ctrl_replacedWayNeedWriteback;
  wire                store_ctrl_refillHit;
  wire                store_ctrl_lineBusy;
  wire                store_ctrl_waysHitHazard;
  wire                store_ctrl_wasClean;
  wire                store_ctrl_bankBusy;
  wire                store_ctrl_hitFault;
  wire       [0:0]    store_ctrl_refillWay;
  wire                store_ctrl_canRefill;
  wire                store_ctrl_askRefill;
  reg                 store_ctrl_startRefill;
  reg                 store_ctrl_writeCache;
  reg                 store_ctrl_setDirty;
  wire                _zz_store_ctrl_wayId;
  wire       [0:0]    store_ctrl_wayId;
  wire       [1:0]    store_ctrl_needFlushs;
  wire       [1:0]    _zz_store_ctrl_needFlushs_bools_0;
  wire                store_ctrl_needFlushs_bools_0;
  wire                store_ctrl_needFlushs_bools_1;
  reg        [1:0]    _zz_store_ctrl_needFlushOh;
  wire       [1:0]    store_ctrl_needFlushOh;
  wire                _zz_store_ctrl_needFlushSel;
  wire       [0:0]    store_ctrl_needFlushSel;
  wire                store_ctrl_needFlush;
  wire                store_ctrl_canFlush;
  wire                store_ctrl_startFlush;
  wire                when_dcache2_l1542;
  wire                when_dcache2_l1552;
  wire                when_dcache2_l1583;
  wire                when_dcache2_l1583_1;
  wire       [31:0]   _zz_39;
  wire       [3:0]    _zz_40;
  wire       [3:0]    _zz_41;
  wire       [0:0]    _zz_42;
  wire       [0:0]    _zz_43;
  wire       [0:0]    _zz_44;
  wire       [0:0]    _zz_45;
  wire       [0:0]    _zz_46;
  wire       [0:0]    _zz_47;
  wire                when_Pipeline_l276_2;
  wire                when_Pipeline_l276_3;
  (* ram_style = "block" *) reg [7:0] banks_0_mem_symbol0 [0:127];
  (* ram_style = "block" *) reg [7:0] banks_0_mem_symbol1 [0:127];
  (* ram_style = "block" *) reg [7:0] banks_0_mem_symbol2 [0:127];
  (* ram_style = "block" *) reg [7:0] banks_0_mem_symbol3 [0:127];
  reg [7:0] _zz_banks_0_memsymbol_read;
  reg [7:0] _zz_banks_0_memsymbol_read_1;
  reg [7:0] _zz_banks_0_memsymbol_read_2;
  reg [7:0] _zz_banks_0_memsymbol_read_3;
  (* ram_style = "block" *) reg [7:0] banks_1_mem_symbol0 [0:127];
  (* ram_style = "block" *) reg [7:0] banks_1_mem_symbol1 [0:127];
  (* ram_style = "block" *) reg [7:0] banks_1_mem_symbol2 [0:127];
  (* ram_style = "block" *) reg [7:0] banks_1_mem_symbol3 [0:127];
  reg [7:0] _zz_banks_1_memsymbol_read;
  reg [7:0] _zz_banks_1_memsymbol_read_1;
  reg [7:0] _zz_banks_1_memsymbol_read_2;
  reg [7:0] _zz_banks_1_memsymbol_read_3;
  (* ram_style = "distributed" *) reg [24:0] ways_0_mem [0:15];
  (* ram_style = "distributed" *) reg [24:0] ways_1_mem [0:15];
  (* ram_style = "distributed" *) reg [1:0] status_mem [0:15];
  (* ram_style = "block" *) reg [31:0] writeback_victimBuffer [0:63];

  assign _zz_status_loadRead_rsp_0_dirty_1 = _zz_status_loadRead_rsp_0_dirty[0 : 0];
  assign _zz_status_loadRead_rsp_1_dirty = _zz_status_loadRead_rsp_0_dirty[1 : 1];
  assign _zz_status_storeRead_rsp_0_dirty_1 = _zz_status_storeRead_rsp_0_dirty[0 : 0];
  assign _zz_status_storeRead_rsp_1_dirty = _zz_status_storeRead_rsp_0_dirty[1 : 1];
  assign _zz__zz_refill_free_1 = (_zz_refill_free - 8'h01);
  assign _zz__zz_writeback_free_1 = (_zz_writeback_free - 8'h01);
  assign _zz_writeback_read_wordIndex_1 = writeback_read_slotRead_valid;
  assign _zz_writeback_read_wordIndex = {2'd0, _zz_writeback_read_wordIndex_1};
  assign _zz_writeback_write_wordIndex_1 = writeback_write_bufferRead_fire;
  assign _zz_writeback_write_wordIndex = {2'd0, _zz_writeback_write_wordIndex_1};
  assign _zz_when = 1'b1;
  assign _zz_when_1 = 1'b1;
  assign _zz_ways_0_mem_port = {waysWrite_tag_fault,{waysWrite_tag_address,waysWrite_tag_loaded}};
  assign _zz_ways_0_mem_port_1 = waysWrite_mask[0];
  assign _zz_ways_1_mem_port = {waysWrite_tag_fault,{waysWrite_tag_address,waysWrite_tag_loaded}};
  assign _zz_ways_1_mem_port_1 = waysWrite_mask[1];
  assign _zz_status_mem_port = {status_write_payload_data_1_dirty,status_write_payload_data_0_dirty};
  assign _zz_writeback_victimBuffer_port = {writeback_read_slotReadLast_payload_id,writeback_read_slotReadLast_payload_wordIndex};
  assign _zz_refill_read_arbiter_oh = refill_read_arbiter_hits[6];
  assign _zz_refill_read_arbiter_oh_1 = refill_read_arbiter_hits[5];
  assign _zz_refill_read_arbiter_oh_2 = {_zz_refill_read_arbiter_oh_3,{_zz_refill_read_arbiter_oh_4,_zz_refill_read_arbiter_oh_5}};
  assign _zz_refill_read_arbiter_oh_9 = refill_read_arbiter_hits[7];
  assign _zz_refill_read_arbiter_oh_10 = {_zz_refill_read_arbiter_oh_11,{_zz_refill_read_arbiter_oh_12,_zz_refill_read_arbiter_oh_13}};
  assign _zz_refill_read_arbiter_oh_19 = {_zz_refill_read_arbiter_oh_20,{_zz_refill_read_arbiter_oh_21,_zz_refill_read_arbiter_oh_22}};
  assign _zz_refill_read_arbiter_oh_29 = ({_zz_refill_read_arbiter_oh_30,_zz_refill_read_arbiter_oh_31} & refill_slots_4_priority);
  assign _zz_refill_read_arbiter_oh_38 = 7'h0;
  assign _zz_refill_read_arbiter_oh_39 = ((_zz_refill_read_arbiter_oh_40 & refill_slots_3_priority) == 7'h0);
  assign _zz_refill_read_arbiter_oh_49 = (_zz_refill_read_arbiter_oh_50 == _zz_refill_read_arbiter_oh_59);
  assign _zz_refill_read_arbiter_oh_60 = {_zz_refill_read_arbiter_oh_61,_zz_refill_read_arbiter_oh_69};
  assign _zz_refill_read_arbiter_oh_3 = refill_read_arbiter_hits[4];
  assign _zz_refill_read_arbiter_oh_4 = refill_read_arbiter_hits[3];
  assign _zz_refill_read_arbiter_oh_5 = {_zz_refill_read_arbiter_oh_6,{_zz_refill_read_arbiter_oh_7,_zz_refill_read_arbiter_oh_8}};
  assign _zz_refill_read_arbiter_oh_11 = refill_read_arbiter_hits[5];
  assign _zz_refill_read_arbiter_oh_12 = refill_read_arbiter_hits[4];
  assign _zz_refill_read_arbiter_oh_13 = {_zz_refill_read_arbiter_oh_14,{_zz_refill_read_arbiter_oh_15,_zz_refill_read_arbiter_oh_16}};
  assign _zz_refill_read_arbiter_oh_20 = refill_read_arbiter_hits[7];
  assign _zz_refill_read_arbiter_oh_21 = refill_read_arbiter_hits[6];
  assign _zz_refill_read_arbiter_oh_22 = {_zz_refill_read_arbiter_oh_23,{_zz_refill_read_arbiter_oh_24,_zz_refill_read_arbiter_oh_25}};
  assign _zz_refill_read_arbiter_oh_30 = refill_read_arbiter_hits[7];
  assign _zz_refill_read_arbiter_oh_31 = {_zz_refill_read_arbiter_oh_32,{_zz_refill_read_arbiter_oh_33,_zz_refill_read_arbiter_oh_34}};
  assign _zz_refill_read_arbiter_oh_40 = {_zz_refill_read_arbiter_oh_41,{_zz_refill_read_arbiter_oh_42,_zz_refill_read_arbiter_oh_43}};
  assign _zz_refill_read_arbiter_oh_50 = ({_zz_refill_read_arbiter_oh_51,_zz_refill_read_arbiter_oh_52} & refill_slots_2_priority);
  assign _zz_refill_read_arbiter_oh_59 = 7'h0;
  assign _zz_refill_read_arbiter_oh_61 = ((_zz_refill_read_arbiter_oh_62 & refill_slots_1_priority) == 7'h0);
  assign _zz_refill_read_arbiter_oh_69 = ((_zz_refill_read_arbiter_oh_70 & refill_slots_0_priority) == 7'h0);
  assign _zz_refill_read_arbiter_oh_6 = refill_read_arbiter_hits[2];
  assign _zz_refill_read_arbiter_oh_7 = refill_read_arbiter_hits[1];
  assign _zz_refill_read_arbiter_oh_8 = refill_read_arbiter_hits[0];
  assign _zz_refill_read_arbiter_oh_14 = refill_read_arbiter_hits[3];
  assign _zz_refill_read_arbiter_oh_15 = refill_read_arbiter_hits[2];
  assign _zz_refill_read_arbiter_oh_16 = {_zz_refill_read_arbiter_oh_17,_zz_refill_read_arbiter_oh_18};
  assign _zz_refill_read_arbiter_oh_23 = refill_read_arbiter_hits[4];
  assign _zz_refill_read_arbiter_oh_24 = refill_read_arbiter_hits[3];
  assign _zz_refill_read_arbiter_oh_25 = {_zz_refill_read_arbiter_oh_26,{_zz_refill_read_arbiter_oh_27,_zz_refill_read_arbiter_oh_28}};
  assign _zz_refill_read_arbiter_oh_32 = refill_read_arbiter_hits[6];
  assign _zz_refill_read_arbiter_oh_33 = refill_read_arbiter_hits[5];
  assign _zz_refill_read_arbiter_oh_34 = {_zz_refill_read_arbiter_oh_35,{_zz_refill_read_arbiter_oh_36,_zz_refill_read_arbiter_oh_37}};
  assign _zz_refill_read_arbiter_oh_41 = refill_read_arbiter_hits[7];
  assign _zz_refill_read_arbiter_oh_42 = refill_read_arbiter_hits[6];
  assign _zz_refill_read_arbiter_oh_43 = {_zz_refill_read_arbiter_oh_44,{_zz_refill_read_arbiter_oh_45,_zz_refill_read_arbiter_oh_46}};
  assign _zz_refill_read_arbiter_oh_51 = refill_read_arbiter_hits[7];
  assign _zz_refill_read_arbiter_oh_52 = {_zz_refill_read_arbiter_oh_53,{_zz_refill_read_arbiter_oh_54,_zz_refill_read_arbiter_oh_55}};
  assign _zz_refill_read_arbiter_oh_62 = {_zz_refill_read_arbiter_oh_63,{_zz_refill_read_arbiter_oh_64,_zz_refill_read_arbiter_oh_65}};
  assign _zz_refill_read_arbiter_oh_70 = {_zz_refill_read_arbiter_oh_71,{_zz_refill_read_arbiter_oh_72,_zz_refill_read_arbiter_oh_73}};
  assign _zz_refill_read_arbiter_oh_17 = refill_read_arbiter_hits[1];
  assign _zz_refill_read_arbiter_oh_18 = refill_read_arbiter_hits[0];
  assign _zz_refill_read_arbiter_oh_26 = refill_read_arbiter_hits[2];
  assign _zz_refill_read_arbiter_oh_27 = refill_read_arbiter_hits[1];
  assign _zz_refill_read_arbiter_oh_28 = refill_read_arbiter_hits[0];
  assign _zz_refill_read_arbiter_oh_35 = refill_read_arbiter_hits[3];
  assign _zz_refill_read_arbiter_oh_36 = refill_read_arbiter_hits[2];
  assign _zz_refill_read_arbiter_oh_37 = {refill_read_arbiter_hits[1],refill_read_arbiter_hits[0]};
  assign _zz_refill_read_arbiter_oh_44 = refill_read_arbiter_hits[5];
  assign _zz_refill_read_arbiter_oh_45 = refill_read_arbiter_hits[4];
  assign _zz_refill_read_arbiter_oh_46 = {refill_read_arbiter_hits[2],{_zz_refill_read_arbiter_oh_47,_zz_refill_read_arbiter_oh_48}};
  assign _zz_refill_read_arbiter_oh_53 = refill_read_arbiter_hits[6];
  assign _zz_refill_read_arbiter_oh_54 = refill_read_arbiter_hits[5];
  assign _zz_refill_read_arbiter_oh_55 = {refill_read_arbiter_hits[4],{_zz_refill_read_arbiter_oh_56,{_zz_refill_read_arbiter_oh_57,_zz_refill_read_arbiter_oh_58}}};
  assign _zz_refill_read_arbiter_oh_63 = refill_read_arbiter_hits[7];
  assign _zz_refill_read_arbiter_oh_64 = refill_read_arbiter_hits[6];
  assign _zz_refill_read_arbiter_oh_65 = {refill_read_arbiter_hits[5],{_zz_refill_read_arbiter_oh_66,{_zz_refill_read_arbiter_oh_67,_zz_refill_read_arbiter_oh_68}}};
  assign _zz_refill_read_arbiter_oh_71 = refill_read_arbiter_hits[7];
  assign _zz_refill_read_arbiter_oh_72 = refill_read_arbiter_hits[6];
  assign _zz_refill_read_arbiter_oh_73 = {refill_read_arbiter_hits[5],{_zz_refill_read_arbiter_oh_74,{_zz_refill_read_arbiter_oh_75,_zz_refill_read_arbiter_oh_76}}};
  assign _zz_refill_read_arbiter_oh_47 = refill_read_arbiter_hits[1];
  assign _zz_refill_read_arbiter_oh_48 = refill_read_arbiter_hits[0];
  assign _zz_refill_read_arbiter_oh_56 = refill_read_arbiter_hits[3];
  assign _zz_refill_read_arbiter_oh_57 = refill_read_arbiter_hits[1];
  assign _zz_refill_read_arbiter_oh_58 = refill_read_arbiter_hits[0];
  assign _zz_refill_read_arbiter_oh_66 = refill_read_arbiter_hits[4];
  assign _zz_refill_read_arbiter_oh_67 = refill_read_arbiter_hits[3];
  assign _zz_refill_read_arbiter_oh_68 = {refill_read_arbiter_hits[2],refill_read_arbiter_hits[0]};
  assign _zz_refill_read_arbiter_oh_74 = refill_read_arbiter_hits[4];
  assign _zz_refill_read_arbiter_oh_75 = refill_read_arbiter_hits[3];
  assign _zz_refill_read_arbiter_oh_76 = {refill_read_arbiter_hits[2],refill_read_arbiter_hits[1]};
  assign _zz_writeback_read_arbiter_oh = writeback_read_arbiter_hits[6];
  assign _zz_writeback_read_arbiter_oh_1 = writeback_read_arbiter_hits[5];
  assign _zz_writeback_read_arbiter_oh_2 = {_zz_writeback_read_arbiter_oh_3,{_zz_writeback_read_arbiter_oh_4,_zz_writeback_read_arbiter_oh_5}};
  assign _zz_writeback_read_arbiter_oh_9 = writeback_read_arbiter_hits[7];
  assign _zz_writeback_read_arbiter_oh_10 = {_zz_writeback_read_arbiter_oh_11,{_zz_writeback_read_arbiter_oh_12,_zz_writeback_read_arbiter_oh_13}};
  assign _zz_writeback_read_arbiter_oh_19 = {_zz_writeback_read_arbiter_oh_20,{_zz_writeback_read_arbiter_oh_21,_zz_writeback_read_arbiter_oh_22}};
  assign _zz_writeback_read_arbiter_oh_29 = ({_zz_writeback_read_arbiter_oh_30,_zz_writeback_read_arbiter_oh_31} & writeback_slots_4_priority);
  assign _zz_writeback_read_arbiter_oh_38 = 7'h0;
  assign _zz_writeback_read_arbiter_oh_39 = ((_zz_writeback_read_arbiter_oh_40 & writeback_slots_3_priority) == 7'h0);
  assign _zz_writeback_read_arbiter_oh_49 = (_zz_writeback_read_arbiter_oh_50 == _zz_writeback_read_arbiter_oh_59);
  assign _zz_writeback_read_arbiter_oh_60 = {_zz_writeback_read_arbiter_oh_61,_zz_writeback_read_arbiter_oh_69};
  assign _zz_writeback_read_arbiter_oh_3 = writeback_read_arbiter_hits[4];
  assign _zz_writeback_read_arbiter_oh_4 = writeback_read_arbiter_hits[3];
  assign _zz_writeback_read_arbiter_oh_5 = {_zz_writeback_read_arbiter_oh_6,{_zz_writeback_read_arbiter_oh_7,_zz_writeback_read_arbiter_oh_8}};
  assign _zz_writeback_read_arbiter_oh_11 = writeback_read_arbiter_hits[5];
  assign _zz_writeback_read_arbiter_oh_12 = writeback_read_arbiter_hits[4];
  assign _zz_writeback_read_arbiter_oh_13 = {_zz_writeback_read_arbiter_oh_14,{_zz_writeback_read_arbiter_oh_15,_zz_writeback_read_arbiter_oh_16}};
  assign _zz_writeback_read_arbiter_oh_20 = writeback_read_arbiter_hits[7];
  assign _zz_writeback_read_arbiter_oh_21 = writeback_read_arbiter_hits[6];
  assign _zz_writeback_read_arbiter_oh_22 = {_zz_writeback_read_arbiter_oh_23,{_zz_writeback_read_arbiter_oh_24,_zz_writeback_read_arbiter_oh_25}};
  assign _zz_writeback_read_arbiter_oh_30 = writeback_read_arbiter_hits[7];
  assign _zz_writeback_read_arbiter_oh_31 = {_zz_writeback_read_arbiter_oh_32,{_zz_writeback_read_arbiter_oh_33,_zz_writeback_read_arbiter_oh_34}};
  assign _zz_writeback_read_arbiter_oh_40 = {_zz_writeback_read_arbiter_oh_41,{_zz_writeback_read_arbiter_oh_42,_zz_writeback_read_arbiter_oh_43}};
  assign _zz_writeback_read_arbiter_oh_50 = ({_zz_writeback_read_arbiter_oh_51,_zz_writeback_read_arbiter_oh_52} & writeback_slots_2_priority);
  assign _zz_writeback_read_arbiter_oh_59 = 7'h0;
  assign _zz_writeback_read_arbiter_oh_61 = ((_zz_writeback_read_arbiter_oh_62 & writeback_slots_1_priority) == 7'h0);
  assign _zz_writeback_read_arbiter_oh_69 = ((_zz_writeback_read_arbiter_oh_70 & writeback_slots_0_priority) == 7'h0);
  assign _zz_writeback_read_arbiter_oh_6 = writeback_read_arbiter_hits[2];
  assign _zz_writeback_read_arbiter_oh_7 = writeback_read_arbiter_hits[1];
  assign _zz_writeback_read_arbiter_oh_8 = writeback_read_arbiter_hits[0];
  assign _zz_writeback_read_arbiter_oh_14 = writeback_read_arbiter_hits[3];
  assign _zz_writeback_read_arbiter_oh_15 = writeback_read_arbiter_hits[2];
  assign _zz_writeback_read_arbiter_oh_16 = {_zz_writeback_read_arbiter_oh_17,_zz_writeback_read_arbiter_oh_18};
  assign _zz_writeback_read_arbiter_oh_23 = writeback_read_arbiter_hits[4];
  assign _zz_writeback_read_arbiter_oh_24 = writeback_read_arbiter_hits[3];
  assign _zz_writeback_read_arbiter_oh_25 = {_zz_writeback_read_arbiter_oh_26,{_zz_writeback_read_arbiter_oh_27,_zz_writeback_read_arbiter_oh_28}};
  assign _zz_writeback_read_arbiter_oh_32 = writeback_read_arbiter_hits[6];
  assign _zz_writeback_read_arbiter_oh_33 = writeback_read_arbiter_hits[5];
  assign _zz_writeback_read_arbiter_oh_34 = {_zz_writeback_read_arbiter_oh_35,{_zz_writeback_read_arbiter_oh_36,_zz_writeback_read_arbiter_oh_37}};
  assign _zz_writeback_read_arbiter_oh_41 = writeback_read_arbiter_hits[7];
  assign _zz_writeback_read_arbiter_oh_42 = writeback_read_arbiter_hits[6];
  assign _zz_writeback_read_arbiter_oh_43 = {_zz_writeback_read_arbiter_oh_44,{_zz_writeback_read_arbiter_oh_45,_zz_writeback_read_arbiter_oh_46}};
  assign _zz_writeback_read_arbiter_oh_51 = writeback_read_arbiter_hits[7];
  assign _zz_writeback_read_arbiter_oh_52 = {_zz_writeback_read_arbiter_oh_53,{_zz_writeback_read_arbiter_oh_54,_zz_writeback_read_arbiter_oh_55}};
  assign _zz_writeback_read_arbiter_oh_62 = {_zz_writeback_read_arbiter_oh_63,{_zz_writeback_read_arbiter_oh_64,_zz_writeback_read_arbiter_oh_65}};
  assign _zz_writeback_read_arbiter_oh_70 = {_zz_writeback_read_arbiter_oh_71,{_zz_writeback_read_arbiter_oh_72,_zz_writeback_read_arbiter_oh_73}};
  assign _zz_writeback_read_arbiter_oh_17 = writeback_read_arbiter_hits[1];
  assign _zz_writeback_read_arbiter_oh_18 = writeback_read_arbiter_hits[0];
  assign _zz_writeback_read_arbiter_oh_26 = writeback_read_arbiter_hits[2];
  assign _zz_writeback_read_arbiter_oh_27 = writeback_read_arbiter_hits[1];
  assign _zz_writeback_read_arbiter_oh_28 = writeback_read_arbiter_hits[0];
  assign _zz_writeback_read_arbiter_oh_35 = writeback_read_arbiter_hits[3];
  assign _zz_writeback_read_arbiter_oh_36 = writeback_read_arbiter_hits[2];
  assign _zz_writeback_read_arbiter_oh_37 = {writeback_read_arbiter_hits[1],writeback_read_arbiter_hits[0]};
  assign _zz_writeback_read_arbiter_oh_44 = writeback_read_arbiter_hits[5];
  assign _zz_writeback_read_arbiter_oh_45 = writeback_read_arbiter_hits[4];
  assign _zz_writeback_read_arbiter_oh_46 = {writeback_read_arbiter_hits[2],{_zz_writeback_read_arbiter_oh_47,_zz_writeback_read_arbiter_oh_48}};
  assign _zz_writeback_read_arbiter_oh_53 = writeback_read_arbiter_hits[6];
  assign _zz_writeback_read_arbiter_oh_54 = writeback_read_arbiter_hits[5];
  assign _zz_writeback_read_arbiter_oh_55 = {writeback_read_arbiter_hits[4],{_zz_writeback_read_arbiter_oh_56,{_zz_writeback_read_arbiter_oh_57,_zz_writeback_read_arbiter_oh_58}}};
  assign _zz_writeback_read_arbiter_oh_63 = writeback_read_arbiter_hits[7];
  assign _zz_writeback_read_arbiter_oh_64 = writeback_read_arbiter_hits[6];
  assign _zz_writeback_read_arbiter_oh_65 = {writeback_read_arbiter_hits[5],{_zz_writeback_read_arbiter_oh_66,{_zz_writeback_read_arbiter_oh_67,_zz_writeback_read_arbiter_oh_68}}};
  assign _zz_writeback_read_arbiter_oh_71 = writeback_read_arbiter_hits[7];
  assign _zz_writeback_read_arbiter_oh_72 = writeback_read_arbiter_hits[6];
  assign _zz_writeback_read_arbiter_oh_73 = {writeback_read_arbiter_hits[5],{_zz_writeback_read_arbiter_oh_74,{_zz_writeback_read_arbiter_oh_75,_zz_writeback_read_arbiter_oh_76}}};
  assign _zz_writeback_read_arbiter_oh_47 = writeback_read_arbiter_hits[1];
  assign _zz_writeback_read_arbiter_oh_48 = writeback_read_arbiter_hits[0];
  assign _zz_writeback_read_arbiter_oh_56 = writeback_read_arbiter_hits[3];
  assign _zz_writeback_read_arbiter_oh_57 = writeback_read_arbiter_hits[1];
  assign _zz_writeback_read_arbiter_oh_58 = writeback_read_arbiter_hits[0];
  assign _zz_writeback_read_arbiter_oh_66 = writeback_read_arbiter_hits[4];
  assign _zz_writeback_read_arbiter_oh_67 = writeback_read_arbiter_hits[3];
  assign _zz_writeback_read_arbiter_oh_68 = {writeback_read_arbiter_hits[2],writeback_read_arbiter_hits[0]};
  assign _zz_writeback_read_arbiter_oh_74 = writeback_read_arbiter_hits[4];
  assign _zz_writeback_read_arbiter_oh_75 = writeback_read_arbiter_hits[3];
  assign _zz_writeback_read_arbiter_oh_76 = {writeback_read_arbiter_hits[2],writeback_read_arbiter_hits[1]};
  assign _zz_writeback_write_arbiter_oh = writeback_write_arbiter_hits[6];
  assign _zz_writeback_write_arbiter_oh_1 = writeback_write_arbiter_hits[5];
  assign _zz_writeback_write_arbiter_oh_2 = {_zz_writeback_write_arbiter_oh_3,{_zz_writeback_write_arbiter_oh_4,_zz_writeback_write_arbiter_oh_5}};
  assign _zz_writeback_write_arbiter_oh_9 = writeback_write_arbiter_hits[7];
  assign _zz_writeback_write_arbiter_oh_10 = {_zz_writeback_write_arbiter_oh_11,{_zz_writeback_write_arbiter_oh_12,_zz_writeback_write_arbiter_oh_13}};
  assign _zz_writeback_write_arbiter_oh_19 = {_zz_writeback_write_arbiter_oh_20,{_zz_writeback_write_arbiter_oh_21,_zz_writeback_write_arbiter_oh_22}};
  assign _zz_writeback_write_arbiter_oh_29 = ({_zz_writeback_write_arbiter_oh_30,_zz_writeback_write_arbiter_oh_31} & writeback_slots_4_priority);
  assign _zz_writeback_write_arbiter_oh_38 = 7'h0;
  assign _zz_writeback_write_arbiter_oh_39 = ((_zz_writeback_write_arbiter_oh_40 & writeback_slots_3_priority) == 7'h0);
  assign _zz_writeback_write_arbiter_oh_49 = (_zz_writeback_write_arbiter_oh_50 == _zz_writeback_write_arbiter_oh_59);
  assign _zz_writeback_write_arbiter_oh_60 = {_zz_writeback_write_arbiter_oh_61,_zz_writeback_write_arbiter_oh_69};
  assign _zz_writeback_write_arbiter_oh_3 = writeback_write_arbiter_hits[4];
  assign _zz_writeback_write_arbiter_oh_4 = writeback_write_arbiter_hits[3];
  assign _zz_writeback_write_arbiter_oh_5 = {_zz_writeback_write_arbiter_oh_6,{_zz_writeback_write_arbiter_oh_7,_zz_writeback_write_arbiter_oh_8}};
  assign _zz_writeback_write_arbiter_oh_11 = writeback_write_arbiter_hits[5];
  assign _zz_writeback_write_arbiter_oh_12 = writeback_write_arbiter_hits[4];
  assign _zz_writeback_write_arbiter_oh_13 = {_zz_writeback_write_arbiter_oh_14,{_zz_writeback_write_arbiter_oh_15,_zz_writeback_write_arbiter_oh_16}};
  assign _zz_writeback_write_arbiter_oh_20 = writeback_write_arbiter_hits[7];
  assign _zz_writeback_write_arbiter_oh_21 = writeback_write_arbiter_hits[6];
  assign _zz_writeback_write_arbiter_oh_22 = {_zz_writeback_write_arbiter_oh_23,{_zz_writeback_write_arbiter_oh_24,_zz_writeback_write_arbiter_oh_25}};
  assign _zz_writeback_write_arbiter_oh_30 = writeback_write_arbiter_hits[7];
  assign _zz_writeback_write_arbiter_oh_31 = {_zz_writeback_write_arbiter_oh_32,{_zz_writeback_write_arbiter_oh_33,_zz_writeback_write_arbiter_oh_34}};
  assign _zz_writeback_write_arbiter_oh_40 = {_zz_writeback_write_arbiter_oh_41,{_zz_writeback_write_arbiter_oh_42,_zz_writeback_write_arbiter_oh_43}};
  assign _zz_writeback_write_arbiter_oh_50 = ({_zz_writeback_write_arbiter_oh_51,_zz_writeback_write_arbiter_oh_52} & writeback_slots_2_priority);
  assign _zz_writeback_write_arbiter_oh_59 = 7'h0;
  assign _zz_writeback_write_arbiter_oh_61 = ((_zz_writeback_write_arbiter_oh_62 & writeback_slots_1_priority) == 7'h0);
  assign _zz_writeback_write_arbiter_oh_69 = ((_zz_writeback_write_arbiter_oh_70 & writeback_slots_0_priority) == 7'h0);
  assign _zz_writeback_write_arbiter_oh_6 = writeback_write_arbiter_hits[2];
  assign _zz_writeback_write_arbiter_oh_7 = writeback_write_arbiter_hits[1];
  assign _zz_writeback_write_arbiter_oh_8 = writeback_write_arbiter_hits[0];
  assign _zz_writeback_write_arbiter_oh_14 = writeback_write_arbiter_hits[3];
  assign _zz_writeback_write_arbiter_oh_15 = writeback_write_arbiter_hits[2];
  assign _zz_writeback_write_arbiter_oh_16 = {_zz_writeback_write_arbiter_oh_17,_zz_writeback_write_arbiter_oh_18};
  assign _zz_writeback_write_arbiter_oh_23 = writeback_write_arbiter_hits[4];
  assign _zz_writeback_write_arbiter_oh_24 = writeback_write_arbiter_hits[3];
  assign _zz_writeback_write_arbiter_oh_25 = {_zz_writeback_write_arbiter_oh_26,{_zz_writeback_write_arbiter_oh_27,_zz_writeback_write_arbiter_oh_28}};
  assign _zz_writeback_write_arbiter_oh_32 = writeback_write_arbiter_hits[6];
  assign _zz_writeback_write_arbiter_oh_33 = writeback_write_arbiter_hits[5];
  assign _zz_writeback_write_arbiter_oh_34 = {_zz_writeback_write_arbiter_oh_35,{_zz_writeback_write_arbiter_oh_36,_zz_writeback_write_arbiter_oh_37}};
  assign _zz_writeback_write_arbiter_oh_41 = writeback_write_arbiter_hits[7];
  assign _zz_writeback_write_arbiter_oh_42 = writeback_write_arbiter_hits[6];
  assign _zz_writeback_write_arbiter_oh_43 = {_zz_writeback_write_arbiter_oh_44,{_zz_writeback_write_arbiter_oh_45,_zz_writeback_write_arbiter_oh_46}};
  assign _zz_writeback_write_arbiter_oh_51 = writeback_write_arbiter_hits[7];
  assign _zz_writeback_write_arbiter_oh_52 = {_zz_writeback_write_arbiter_oh_53,{_zz_writeback_write_arbiter_oh_54,_zz_writeback_write_arbiter_oh_55}};
  assign _zz_writeback_write_arbiter_oh_62 = {_zz_writeback_write_arbiter_oh_63,{_zz_writeback_write_arbiter_oh_64,_zz_writeback_write_arbiter_oh_65}};
  assign _zz_writeback_write_arbiter_oh_70 = {_zz_writeback_write_arbiter_oh_71,{_zz_writeback_write_arbiter_oh_72,_zz_writeback_write_arbiter_oh_73}};
  assign _zz_writeback_write_arbiter_oh_17 = writeback_write_arbiter_hits[1];
  assign _zz_writeback_write_arbiter_oh_18 = writeback_write_arbiter_hits[0];
  assign _zz_writeback_write_arbiter_oh_26 = writeback_write_arbiter_hits[2];
  assign _zz_writeback_write_arbiter_oh_27 = writeback_write_arbiter_hits[1];
  assign _zz_writeback_write_arbiter_oh_28 = writeback_write_arbiter_hits[0];
  assign _zz_writeback_write_arbiter_oh_35 = writeback_write_arbiter_hits[3];
  assign _zz_writeback_write_arbiter_oh_36 = writeback_write_arbiter_hits[2];
  assign _zz_writeback_write_arbiter_oh_37 = {writeback_write_arbiter_hits[1],writeback_write_arbiter_hits[0]};
  assign _zz_writeback_write_arbiter_oh_44 = writeback_write_arbiter_hits[5];
  assign _zz_writeback_write_arbiter_oh_45 = writeback_write_arbiter_hits[4];
  assign _zz_writeback_write_arbiter_oh_46 = {writeback_write_arbiter_hits[2],{_zz_writeback_write_arbiter_oh_47,_zz_writeback_write_arbiter_oh_48}};
  assign _zz_writeback_write_arbiter_oh_53 = writeback_write_arbiter_hits[6];
  assign _zz_writeback_write_arbiter_oh_54 = writeback_write_arbiter_hits[5];
  assign _zz_writeback_write_arbiter_oh_55 = {writeback_write_arbiter_hits[4],{_zz_writeback_write_arbiter_oh_56,{_zz_writeback_write_arbiter_oh_57,_zz_writeback_write_arbiter_oh_58}}};
  assign _zz_writeback_write_arbiter_oh_63 = writeback_write_arbiter_hits[7];
  assign _zz_writeback_write_arbiter_oh_64 = writeback_write_arbiter_hits[6];
  assign _zz_writeback_write_arbiter_oh_65 = {writeback_write_arbiter_hits[5],{_zz_writeback_write_arbiter_oh_66,{_zz_writeback_write_arbiter_oh_67,_zz_writeback_write_arbiter_oh_68}}};
  assign _zz_writeback_write_arbiter_oh_71 = writeback_write_arbiter_hits[7];
  assign _zz_writeback_write_arbiter_oh_72 = writeback_write_arbiter_hits[6];
  assign _zz_writeback_write_arbiter_oh_73 = {writeback_write_arbiter_hits[5],{_zz_writeback_write_arbiter_oh_74,{_zz_writeback_write_arbiter_oh_75,_zz_writeback_write_arbiter_oh_76}}};
  assign _zz_writeback_write_arbiter_oh_47 = writeback_write_arbiter_hits[1];
  assign _zz_writeback_write_arbiter_oh_48 = writeback_write_arbiter_hits[0];
  assign _zz_writeback_write_arbiter_oh_56 = writeback_write_arbiter_hits[3];
  assign _zz_writeback_write_arbiter_oh_57 = writeback_write_arbiter_hits[1];
  assign _zz_writeback_write_arbiter_oh_58 = writeback_write_arbiter_hits[0];
  assign _zz_writeback_write_arbiter_oh_66 = writeback_write_arbiter_hits[4];
  assign _zz_writeback_write_arbiter_oh_67 = writeback_write_arbiter_hits[3];
  assign _zz_writeback_write_arbiter_oh_68 = {writeback_write_arbiter_hits[2],writeback_write_arbiter_hits[0]};
  assign _zz_writeback_write_arbiter_oh_74 = writeback_write_arbiter_hits[4];
  assign _zz_writeback_write_arbiter_oh_75 = writeback_write_arbiter_hits[3];
  assign _zz_writeback_write_arbiter_oh_76 = {writeback_write_arbiter_hits[2],writeback_write_arbiter_hits[1]};
  assign _zz_load_pipeline_stages_1_REFILL_HITS_EARLY = refill_slots_5_address[31 : 5];
  assign _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_1 = load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5];
  assign _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_2 = (refill_slots_4_address[31 : 5] == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]);
  assign _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_3 = (refill_slots_3_valid && (refill_slots_3_address[31 : 5] == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]));
  assign _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_4 = (refill_slots_2_valid && (refill_slots_2_address[31 : 5] == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]));
  assign _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_5 = {(refill_slots_1_valid && (refill_slots_1_address[31 : 5] == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5])),(refill_slots_0_valid && (refill_slots_0_address[31 : 5] == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]))};
  assign _zz_load_ctrl_lineBusy = refill_slots_7_address[8 : 5];
  assign _zz_load_ctrl_lineBusy_1 = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_load_ctrl_lineBusy_2 = (refill_slots_6_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_load_ctrl_lineBusy_3 = (refill_slots_5_valid && (_zz_load_ctrl_lineBusy_4 == _zz_load_ctrl_lineBusy_5));
  assign _zz_load_ctrl_lineBusy_6 = (refill_slots_4_valid && _zz_load_ctrl_lineBusy_7);
  assign _zz_load_ctrl_lineBusy_8 = {_zz_load_ctrl_lineBusy_9,{_zz_load_ctrl_lineBusy_10,_zz_load_ctrl_lineBusy_13}};
  assign _zz_load_ctrl_lineBusy_16 = writeback_slots_7_address[8 : 5];
  assign _zz_load_ctrl_lineBusy_17 = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_load_ctrl_lineBusy_18 = (writeback_slots_6_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_load_ctrl_lineBusy_19 = (writeback_slots_5_valid && (_zz_load_ctrl_lineBusy_20 == _zz_load_ctrl_lineBusy_21));
  assign _zz_load_ctrl_lineBusy_22 = (writeback_slots_4_valid && _zz_load_ctrl_lineBusy_23);
  assign _zz_load_ctrl_lineBusy_24 = {_zz_load_ctrl_lineBusy_25,{_zz_load_ctrl_lineBusy_26,_zz_load_ctrl_lineBusy_29}};
  assign _zz_load_ctrl_lineBusy_4 = refill_slots_5_address[8 : 5];
  assign _zz_load_ctrl_lineBusy_5 = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_load_ctrl_lineBusy_7 = (refill_slots_4_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_load_ctrl_lineBusy_9 = (refill_slots_3_valid && (refill_slots_3_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]));
  assign _zz_load_ctrl_lineBusy_10 = (refill_slots_2_valid && (_zz_load_ctrl_lineBusy_11 == _zz_load_ctrl_lineBusy_12));
  assign _zz_load_ctrl_lineBusy_13 = {(refill_slots_1_valid && _zz_load_ctrl_lineBusy_14),(refill_slots_0_valid && _zz_load_ctrl_lineBusy_15)};
  assign _zz_load_ctrl_lineBusy_20 = writeback_slots_5_address[8 : 5];
  assign _zz_load_ctrl_lineBusy_21 = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_load_ctrl_lineBusy_23 = (writeback_slots_4_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_load_ctrl_lineBusy_25 = (writeback_slots_3_valid && (writeback_slots_3_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]));
  assign _zz_load_ctrl_lineBusy_26 = (writeback_slots_2_valid && (_zz_load_ctrl_lineBusy_27 == _zz_load_ctrl_lineBusy_28));
  assign _zz_load_ctrl_lineBusy_29 = {(writeback_slots_1_valid && _zz_load_ctrl_lineBusy_30),(writeback_slots_0_valid && _zz_load_ctrl_lineBusy_31)};
  assign _zz_load_ctrl_lineBusy_11 = refill_slots_2_address[8 : 5];
  assign _zz_load_ctrl_lineBusy_12 = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_load_ctrl_lineBusy_14 = (refill_slots_1_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_load_ctrl_lineBusy_15 = (refill_slots_0_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_load_ctrl_lineBusy_27 = writeback_slots_2_address[8 : 5];
  assign _zz_load_ctrl_lineBusy_28 = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_load_ctrl_lineBusy_30 = (writeback_slots_1_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_load_ctrl_lineBusy_31 = (writeback_slots_0_address[8 : 5] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_store_pipeline_stages_1_REFILL_HITS_EARLY = refill_slots_5_address[31 : 5];
  assign _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_1 = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5];
  assign _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_2 = (refill_slots_4_address[31 : 5] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]);
  assign _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_3 = (refill_slots_3_valid && (refill_slots_3_address[31 : 5] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]));
  assign _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_4 = (refill_slots_2_valid && (refill_slots_2_address[31 : 5] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]));
  assign _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_5 = {(refill_slots_1_valid && (refill_slots_1_address[31 : 5] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5])),(refill_slots_0_valid && (refill_slots_0_address[31 : 5] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]))};
  assign _zz_store_ctrl_lineBusy = refill_slots_7_address[8 : 5];
  assign _zz_store_ctrl_lineBusy_1 = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_store_ctrl_lineBusy_2 = (refill_slots_6_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_store_ctrl_lineBusy_3 = (refill_slots_5_valid && (_zz_store_ctrl_lineBusy_4 == _zz_store_ctrl_lineBusy_5));
  assign _zz_store_ctrl_lineBusy_6 = (refill_slots_4_valid && _zz_store_ctrl_lineBusy_7);
  assign _zz_store_ctrl_lineBusy_8 = {_zz_store_ctrl_lineBusy_9,{_zz_store_ctrl_lineBusy_10,_zz_store_ctrl_lineBusy_13}};
  assign _zz_store_ctrl_lineBusy_16 = writeback_slots_7_address[8 : 5];
  assign _zz_store_ctrl_lineBusy_17 = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_store_ctrl_lineBusy_18 = (writeback_slots_6_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_store_ctrl_lineBusy_19 = (writeback_slots_5_valid && (_zz_store_ctrl_lineBusy_20 == _zz_store_ctrl_lineBusy_21));
  assign _zz_store_ctrl_lineBusy_22 = (writeback_slots_4_valid && _zz_store_ctrl_lineBusy_23);
  assign _zz_store_ctrl_lineBusy_24 = {_zz_store_ctrl_lineBusy_25,{_zz_store_ctrl_lineBusy_26,_zz_store_ctrl_lineBusy_29}};
  assign _zz_store_ctrl_lineBusy_4 = refill_slots_5_address[8 : 5];
  assign _zz_store_ctrl_lineBusy_5 = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_store_ctrl_lineBusy_7 = (refill_slots_4_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_store_ctrl_lineBusy_9 = (refill_slots_3_valid && (refill_slots_3_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]));
  assign _zz_store_ctrl_lineBusy_10 = (refill_slots_2_valid && (_zz_store_ctrl_lineBusy_11 == _zz_store_ctrl_lineBusy_12));
  assign _zz_store_ctrl_lineBusy_13 = {(refill_slots_1_valid && _zz_store_ctrl_lineBusy_14),(refill_slots_0_valid && _zz_store_ctrl_lineBusy_15)};
  assign _zz_store_ctrl_lineBusy_20 = writeback_slots_5_address[8 : 5];
  assign _zz_store_ctrl_lineBusy_21 = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_store_ctrl_lineBusy_23 = (writeback_slots_4_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_store_ctrl_lineBusy_25 = (writeback_slots_3_valid && (writeback_slots_3_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]));
  assign _zz_store_ctrl_lineBusy_26 = (writeback_slots_2_valid && (_zz_store_ctrl_lineBusy_27 == _zz_store_ctrl_lineBusy_28));
  assign _zz_store_ctrl_lineBusy_29 = {(writeback_slots_1_valid && _zz_store_ctrl_lineBusy_30),(writeback_slots_0_valid && _zz_store_ctrl_lineBusy_31)};
  assign _zz_store_ctrl_lineBusy_11 = refill_slots_2_address[8 : 5];
  assign _zz_store_ctrl_lineBusy_12 = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_store_ctrl_lineBusy_14 = (refill_slots_1_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_store_ctrl_lineBusy_15 = (refill_slots_0_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_store_ctrl_lineBusy_27 = writeback_slots_2_address[8 : 5];
  assign _zz_store_ctrl_lineBusy_28 = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_store_ctrl_lineBusy_30 = (writeback_slots_1_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  assign _zz_store_ctrl_lineBusy_31 = (writeback_slots_0_address[8 : 5] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]);
  always @(*) begin
    banks_0_mem_spinal_port1 = {_zz_banks_0_memsymbol_read_3, _zz_banks_0_memsymbol_read_2, _zz_banks_0_memsymbol_read_1, _zz_banks_0_memsymbol_read};
  end
  always @(posedge clk) begin
    if(banks_0_write_payload_mask[0] && banks_0_write_valid) begin
      banks_0_mem_symbol0[banks_0_write_payload_address] <= banks_0_write_payload_data[7 : 0];
    end
    if(banks_0_write_payload_mask[1] && banks_0_write_valid) begin
      banks_0_mem_symbol1[banks_0_write_payload_address] <= banks_0_write_payload_data[15 : 8];
    end
    if(banks_0_write_payload_mask[2] && banks_0_write_valid) begin
      banks_0_mem_symbol2[banks_0_write_payload_address] <= banks_0_write_payload_data[23 : 16];
    end
    if(banks_0_write_payload_mask[3] && banks_0_write_valid) begin
      banks_0_mem_symbol3[banks_0_write_payload_address] <= banks_0_write_payload_data[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(banks_0_read_cmd_valid) begin
      _zz_banks_0_memsymbol_read <= banks_0_mem_symbol0[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_1 <= banks_0_mem_symbol1[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_2 <= banks_0_mem_symbol2[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_3 <= banks_0_mem_symbol3[banks_0_read_cmd_payload];
    end
  end

  always @(*) begin
    banks_1_mem_spinal_port1 = {_zz_banks_1_memsymbol_read_3, _zz_banks_1_memsymbol_read_2, _zz_banks_1_memsymbol_read_1, _zz_banks_1_memsymbol_read};
  end
  always @(posedge clk) begin
    if(banks_1_write_payload_mask[0] && banks_1_write_valid) begin
      banks_1_mem_symbol0[banks_1_write_payload_address] <= banks_1_write_payload_data[7 : 0];
    end
    if(banks_1_write_payload_mask[1] && banks_1_write_valid) begin
      banks_1_mem_symbol1[banks_1_write_payload_address] <= banks_1_write_payload_data[15 : 8];
    end
    if(banks_1_write_payload_mask[2] && banks_1_write_valid) begin
      banks_1_mem_symbol2[banks_1_write_payload_address] <= banks_1_write_payload_data[23 : 16];
    end
    if(banks_1_write_payload_mask[3] && banks_1_write_valid) begin
      banks_1_mem_symbol3[banks_1_write_payload_address] <= banks_1_write_payload_data[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(banks_1_read_cmd_valid) begin
      _zz_banks_1_memsymbol_read <= banks_1_mem_symbol0[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_1 <= banks_1_mem_symbol1[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_2 <= banks_1_mem_symbol2[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_3 <= banks_1_mem_symbol3[banks_1_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_ways_0_mem_port_1) begin
      ways_0_mem[waysWrite_address] <= _zz_ways_0_mem_port;
    end
  end

  assign ways_0_mem_spinal_port1 = ways_0_mem[ways_0_loadRead_cmd_payload];
  assign ways_0_mem_spinal_port2 = ways_0_mem[ways_0_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_ways_1_mem_port_1) begin
      ways_1_mem[waysWrite_address] <= _zz_ways_1_mem_port;
    end
  end

  assign ways_1_mem_spinal_port1 = ways_1_mem[ways_1_loadRead_cmd_payload];
  assign ways_1_mem_spinal_port2 = ways_1_mem[ways_1_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_2) begin
      status_mem[status_write_payload_address] <= _zz_status_mem_port;
    end
  end

  assign status_mem_spinal_port1 = status_mem[status_loadRead_cmd_payload];
  assign status_mem_spinal_port2 = status_mem[status_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_1) begin
      writeback_victimBuffer[_zz_writeback_victimBuffer_port] <= writeback_read_readedData;
    end
  end

  always @(posedge clk) begin
    if(writeback_write_bufferRead_ready) begin
      writeback_victimBuffer_spinal_port1 <= writeback_victimBuffer[_zz_writeback_write_word];
    end
  end

  always @(*) begin
    case(refill_read_arbiter_sel)
      3'b000 : _zz_refill_read_cmdAddress = refill_slots_0_address[31 : 5];
      3'b001 : _zz_refill_read_cmdAddress = refill_slots_1_address[31 : 5];
      3'b010 : _zz_refill_read_cmdAddress = refill_slots_2_address[31 : 5];
      3'b011 : _zz_refill_read_cmdAddress = refill_slots_3_address[31 : 5];
      3'b100 : _zz_refill_read_cmdAddress = refill_slots_4_address[31 : 5];
      3'b101 : _zz_refill_read_cmdAddress = refill_slots_5_address[31 : 5];
      3'b110 : _zz_refill_read_cmdAddress = refill_slots_6_address[31 : 5];
      default : _zz_refill_read_cmdAddress = refill_slots_7_address[31 : 5];
    endcase
  end

  always @(*) begin
    case(io_mem_read_rsp_payload_id)
      3'b000 : begin
        _zz_refill_read_rspAddress = refill_slots_0_address;
        _zz_refill_read_way = refill_slots_0_way;
      end
      3'b001 : begin
        _zz_refill_read_rspAddress = refill_slots_1_address;
        _zz_refill_read_way = refill_slots_1_way;
      end
      3'b010 : begin
        _zz_refill_read_rspAddress = refill_slots_2_address;
        _zz_refill_read_way = refill_slots_2_way;
      end
      3'b011 : begin
        _zz_refill_read_rspAddress = refill_slots_3_address;
        _zz_refill_read_way = refill_slots_3_way;
      end
      3'b100 : begin
        _zz_refill_read_rspAddress = refill_slots_4_address;
        _zz_refill_read_way = refill_slots_4_way;
      end
      3'b101 : begin
        _zz_refill_read_rspAddress = refill_slots_5_address;
        _zz_refill_read_way = refill_slots_5_way;
      end
      3'b110 : begin
        _zz_refill_read_rspAddress = refill_slots_6_address;
        _zz_refill_read_way = refill_slots_6_way;
      end
      default : begin
        _zz_refill_read_rspAddress = refill_slots_7_address;
        _zz_refill_read_way = refill_slots_7_way;
      end
    endcase
  end

  always @(*) begin
    case(writeback_read_arbiter_sel)
      3'b000 : begin
        _zz_writeback_read_address = writeback_slots_0_address;
        _zz_writeback_read_way = writeback_slots_0_way;
      end
      3'b001 : begin
        _zz_writeback_read_address = writeback_slots_1_address;
        _zz_writeback_read_way = writeback_slots_1_way;
      end
      3'b010 : begin
        _zz_writeback_read_address = writeback_slots_2_address;
        _zz_writeback_read_way = writeback_slots_2_way;
      end
      3'b011 : begin
        _zz_writeback_read_address = writeback_slots_3_address;
        _zz_writeback_read_way = writeback_slots_3_way;
      end
      3'b100 : begin
        _zz_writeback_read_address = writeback_slots_4_address;
        _zz_writeback_read_way = writeback_slots_4_way;
      end
      3'b101 : begin
        _zz_writeback_read_address = writeback_slots_5_address;
        _zz_writeback_read_way = writeback_slots_5_way;
      end
      3'b110 : begin
        _zz_writeback_read_address = writeback_slots_6_address;
        _zz_writeback_read_way = writeback_slots_6_way;
      end
      default : begin
        _zz_writeback_read_address = writeback_slots_7_address;
        _zz_writeback_read_way = writeback_slots_7_way;
      end
    endcase
  end

  always @(*) begin
    case(writeback_read_slotReadLast_payload_way)
      1'b0 : _zz_writeback_read_readedData = banks_0_read_rsp;
      default : _zz_writeback_read_readedData = banks_1_read_rsp;
    endcase
  end

  always @(*) begin
    case(writeback_write_arbiter_sel)
      3'b000 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_0_address;
      3'b001 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_1_address;
      3'b010 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_2_address;
      3'b011 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_3_address;
      3'b100 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_4_address;
      3'b101 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_5_address;
      3'b110 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_6_address;
      default : _zz_writeback_write_bufferRead_payload_address = writeback_slots_7_address;
    endcase
  end

  always @(*) begin
    case(load_ctrl_refillWay)
      1'b0 : begin
        _zz__zz_refill_push_payload_victim = load_pipeline_stages_2_STATUS_0_dirty;
        _zz_load_ctrl_refillWayNeedWriteback = load_pipeline_stages_2_WAYS_TAGS_0_loaded;
        _zz_writeback_push_payload_address = load_pipeline_stages_2_WAYS_TAGS_0_address;
      end
      default : begin
        _zz__zz_refill_push_payload_victim = load_pipeline_stages_2_STATUS_1_dirty;
        _zz_load_ctrl_refillWayNeedWriteback = load_pipeline_stages_2_WAYS_TAGS_1_loaded;
        _zz_writeback_push_payload_address = load_pipeline_stages_2_WAYS_TAGS_1_address;
      end
    endcase
  end

  always @(*) begin
    case(store_ctrl_replacedWay)
      1'b0 : begin
        _zz_store_ctrl_replacedWayNeedWriteback = store_pipeline_stages_2_WAYS_TAGS_0_loaded;
        _zz_store_ctrl_replacedWayNeedWriteback_1 = store_pipeline_stages_2_STATUS_0_dirty;
      end
      default : begin
        _zz_store_ctrl_replacedWayNeedWriteback = store_pipeline_stages_2_WAYS_TAGS_1_loaded;
        _zz_store_ctrl_replacedWayNeedWriteback_1 = store_pipeline_stages_2_STATUS_1_dirty;
      end
    endcase
  end

  always @(*) begin
    case(writeback_push_payload_way)
      1'b0 : _zz_writeback_push_payload_address_1 = store_pipeline_stages_2_WAYS_TAGS_0_address;
      default : _zz_writeback_push_payload_address_1 = store_pipeline_stages_2_WAYS_TAGS_1_address;
    endcase
  end

  always @(*) begin
    case(store_ctrl_refillWay)
      1'b0 : _zz_refill_push_payload_victim_1 = store_pipeline_stages_2_STATUS_0_dirty;
      default : _zz_refill_push_payload_victim_1 = store_pipeline_stages_2_STATUS_1_dirty;
    endcase
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(writeback_read_slotReadLast_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(status_write_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    banks_0_read_usedByWriteBack = 1'b0;
    if(when_dcache2_l948) begin
      banks_0_read_usedByWriteBack = 1'b1;
    end
  end

  assign banks_0_read_rsp = banks_0_mem_spinal_port1;
  always @(*) begin
    banks_0_read_cmd_valid = 1'b0;
    if(when_dcache2_l948) begin
      banks_0_read_cmd_valid = 1'b1;
    end
    if(when_dcache2_l1108) begin
      banks_0_read_cmd_valid = (! (load_pipeline_stages_0_valid && (! load_pipeline_stages_0_ready)));
    end
  end

  always @(*) begin
    banks_0_read_cmd_payload = 7'bxxxxxxx;
    if(when_dcache2_l948) begin
      banks_0_read_cmd_payload = {writeback_read_address[8 : 5],writeback_read_wordIndex};
    end
    if(when_dcache2_l1108) begin
      banks_0_read_cmd_payload = load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION[8 : 2];
    end
  end

  always @(*) begin
    banks_1_read_usedByWriteBack = 1'b0;
    if(when_dcache2_l948_1) begin
      banks_1_read_usedByWriteBack = 1'b1;
    end
  end

  assign banks_1_read_rsp = banks_1_mem_spinal_port1;
  always @(*) begin
    banks_1_read_cmd_valid = 1'b0;
    if(when_dcache2_l948_1) begin
      banks_1_read_cmd_valid = 1'b1;
    end
    if(when_dcache2_l1108_1) begin
      banks_1_read_cmd_valid = (! (load_pipeline_stages_0_valid && (! load_pipeline_stages_0_ready)));
    end
  end

  always @(*) begin
    banks_1_read_cmd_payload = 7'bxxxxxxx;
    if(when_dcache2_l948_1) begin
      banks_1_read_cmd_payload = {writeback_read_address[8 : 5],writeback_read_wordIndex};
    end
    if(when_dcache2_l1108_1) begin
      banks_1_read_cmd_payload = load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION[8 : 2];
    end
  end

  always @(*) begin
    waysWrite_mask = 2'b00;
    if(when_dcache2_l680) begin
      waysWrite_mask = 2'b11;
    end
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        waysWrite_mask[refill_read_way] = 1'b1;
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_mask[load_ctrl_refillWay] = 1'b1;
    end
    if(store_ctrl_startRefill) begin
      waysWrite_mask[store_ctrl_refillWay] = 1'b1;
    end
    if(store_ctrl_startFlush) begin
      if(store_pipeline_stages_2_FLUSH_FREE) begin
        if(store_ctrl_needFlushOh[0]) begin
          waysWrite_mask[0] = 1'b1;
        end
        if(_zz_store_ctrl_needFlushSel) begin
          waysWrite_mask[1] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    waysWrite_address = 4'bxxxx;
    if(when_dcache2_l680) begin
      waysWrite_address = invalidate_counter[3:0];
    end
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        waysWrite_address = refill_read_rspAddress[8 : 5];
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_address = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
    end
    if(store_ctrl_startRefill) begin
      waysWrite_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
    end
    if(store_ctrl_startFlush) begin
      if(store_pipeline_stages_2_FLUSH_FREE) begin
        waysWrite_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
      end
    end
  end

  always @(*) begin
    waysWrite_tag_loaded = 1'bx;
    if(when_dcache2_l680) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        waysWrite_tag_loaded = 1'b1;
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(store_ctrl_startRefill) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(store_ctrl_startFlush) begin
      if(store_pipeline_stages_2_FLUSH_FREE) begin
        waysWrite_tag_loaded = 1'b0;
      end
    end
  end

  always @(*) begin
    waysWrite_tag_address = 23'bxxxxxxxxxxxxxxxxxxxxxxx;
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        waysWrite_tag_address = refill_read_rspAddress[31 : 9];
      end
    end
  end

  always @(*) begin
    waysWrite_tag_fault = 1'bx;
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        waysWrite_tag_fault = refill_read_faulty;
      end
    end
  end

  assign _zz_ways_0_loadRead_rsp_loaded = ways_0_mem_spinal_port1;
  assign ways_0_loadRead_rsp_loaded = _zz_ways_0_loadRead_rsp_loaded[0];
  assign ways_0_loadRead_rsp_address = _zz_ways_0_loadRead_rsp_loaded[23 : 1];
  assign ways_0_loadRead_rsp_fault = _zz_ways_0_loadRead_rsp_loaded[24];
  assign _zz_ways_0_storeRead_rsp_loaded = ways_0_mem_spinal_port2;
  assign ways_0_storeRead_rsp_loaded = _zz_ways_0_storeRead_rsp_loaded[0];
  assign ways_0_storeRead_rsp_address = _zz_ways_0_storeRead_rsp_loaded[23 : 1];
  assign ways_0_storeRead_rsp_fault = _zz_ways_0_storeRead_rsp_loaded[24];
  assign _zz_ways_1_loadRead_rsp_loaded = ways_1_mem_spinal_port1;
  assign ways_1_loadRead_rsp_loaded = _zz_ways_1_loadRead_rsp_loaded[0];
  assign ways_1_loadRead_rsp_address = _zz_ways_1_loadRead_rsp_loaded[23 : 1];
  assign ways_1_loadRead_rsp_fault = _zz_ways_1_loadRead_rsp_loaded[24];
  assign _zz_ways_1_storeRead_rsp_loaded = ways_1_mem_spinal_port2;
  assign ways_1_storeRead_rsp_loaded = _zz_ways_1_storeRead_rsp_loaded[0];
  assign ways_1_storeRead_rsp_address = _zz_ways_1_storeRead_rsp_loaded[23 : 1];
  assign ways_1_storeRead_rsp_fault = _zz_ways_1_storeRead_rsp_loaded[24];
  always @(*) begin
    status_write_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      status_write_valid = 1'b1;
    end
    if(when_dcache2_l1542) begin
      status_write_valid = 1'b1;
    end
  end

  always @(*) begin
    status_write_payload_address = 4'bxxxx;
    if(load_ctrl_startRefill) begin
      status_write_payload_address = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
    end
    if(when_dcache2_l1542) begin
      status_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
    end
  end

  always @(*) begin
    status_write_payload_data_0_dirty = 1'bx;
    if(load_ctrl_startRefill) begin
      status_write_payload_data_0_dirty = load_pipeline_stages_2_STATUS_0_dirty;
      if(_zz_34[0]) begin
        status_write_payload_data_0_dirty = 1'b0;
      end
    end
    if(when_dcache2_l1542) begin
      status_write_payload_data_0_dirty = store_pipeline_stages_2_STATUS_0_dirty;
    end
    if(when_dcache2_l1552) begin
      if(store_ctrl_startFlush) begin
        case(store_ctrl_needFlushSel)
          1'b0 : begin
            status_write_payload_data_0_dirty = 1'b0;
          end
          default : begin
          end
        endcase
      end
    end
    if(store_ctrl_startRefill) begin
      case(store_ctrl_refillWay)
        1'b0 : begin
          status_write_payload_data_0_dirty = 1'b0;
        end
        default : begin
        end
      endcase
    end
    if(store_ctrl_setDirty) begin
      if(store_pipeline_stages_2_WAYS_HITS[0]) begin
        status_write_payload_data_0_dirty = 1'b1;
      end
    end
  end

  always @(*) begin
    status_write_payload_data_1_dirty = 1'bx;
    if(load_ctrl_startRefill) begin
      status_write_payload_data_1_dirty = load_pipeline_stages_2_STATUS_1_dirty;
      if(_zz_34[1]) begin
        status_write_payload_data_1_dirty = 1'b0;
      end
    end
    if(when_dcache2_l1542) begin
      status_write_payload_data_1_dirty = store_pipeline_stages_2_STATUS_1_dirty;
    end
    if(when_dcache2_l1552) begin
      if(store_ctrl_startFlush) begin
        case(store_ctrl_needFlushSel)
          1'b0 : begin
          end
          default : begin
            status_write_payload_data_1_dirty = 1'b0;
          end
        endcase
      end
    end
    if(store_ctrl_startRefill) begin
      case(store_ctrl_refillWay)
        1'b0 : begin
        end
        default : begin
          status_write_payload_data_1_dirty = 1'b0;
        end
      endcase
    end
    if(store_ctrl_setDirty) begin
      if(_zz_store_ctrl_wayId) begin
        status_write_payload_data_1_dirty = 1'b1;
      end
    end
  end

  assign _zz_status_loadRead_rsp_0_dirty = status_mem_spinal_port1;
  assign status_loadRead_rsp_0_dirty = _zz_status_loadRead_rsp_0_dirty_1[0];
  assign status_loadRead_rsp_1_dirty = _zz_status_loadRead_rsp_1_dirty[0];
  assign _zz_status_storeRead_rsp_0_dirty = status_mem_spinal_port2;
  assign status_storeRead_rsp_0_dirty = _zz_status_storeRead_rsp_0_dirty_1[0];
  assign status_storeRead_rsp_1_dirty = _zz_status_storeRead_rsp_1_dirty[0];
  assign wayRandom_willClear = 1'b0;
  assign wayRandom_willOverflowIfInc = (wayRandom_value == 1'b1);
  assign wayRandom_willOverflow = (wayRandom_willOverflowIfInc && wayRandom_willIncrement);
  always @(*) begin
    wayRandom_valueNext = (wayRandom_value + wayRandom_willIncrement);
    if(wayRandom_willClear) begin
      wayRandom_valueNext = 1'b0;
    end
  end

  assign wayRandom_willIncrement = 1'b1;
  assign invalidate_done = invalidate_counter[4];
  always @(*) begin
    invalidate_reservation_take = 1'b0;
    if(when_dcache2_l680) begin
      invalidate_reservation_take = 1'b1;
    end
  end

  assign when_dcache2_l680 = ((! invalidate_done) && invalidate_reservation_win);
  assign refill_slots_0_loadedDone = (refill_slots_0_loadedCounter == 1'b1);
  assign refill_slots_0_free = (! refill_slots_0_valid);
  assign refill_slots_1_loadedDone = (refill_slots_1_loadedCounter == 1'b1);
  assign refill_slots_1_free = (! refill_slots_1_valid);
  assign refill_slots_2_loadedDone = (refill_slots_2_loadedCounter == 1'b1);
  assign refill_slots_2_free = (! refill_slots_2_valid);
  assign refill_slots_3_loadedDone = (refill_slots_3_loadedCounter == 1'b1);
  assign refill_slots_3_free = (! refill_slots_3_valid);
  assign refill_slots_4_loadedDone = (refill_slots_4_loadedCounter == 1'b1);
  assign refill_slots_4_free = (! refill_slots_4_valid);
  assign refill_slots_5_loadedDone = (refill_slots_5_loadedCounter == 1'b1);
  assign refill_slots_5_free = (! refill_slots_5_valid);
  assign refill_slots_6_loadedDone = (refill_slots_6_loadedCounter == 1'b1);
  assign refill_slots_6_free = (! refill_slots_6_valid);
  assign refill_slots_7_loadedDone = (refill_slots_7_loadedCounter == 1'b1);
  assign refill_slots_7_free = (! refill_slots_7_valid);
  assign _zz_refill_free = {refill_slots_7_free,{refill_slots_6_free,{refill_slots_5_free,{refill_slots_4_free,{refill_slots_3_free,{refill_slots_2_free,{refill_slots_1_free,refill_slots_0_free}}}}}}};
  assign _zz_refill_free_1 = (_zz_refill_free & (~ _zz__zz_refill_free_1));
  assign refill_free = {_zz_refill_free_1[7],{_zz_refill_free_1[6],{_zz_refill_free_1[5],{_zz_refill_free_1[4],{_zz_refill_free_1[3],{_zz_refill_free_1[2],{_zz_refill_free_1[1],refill_slots_0_free}}}}}}};
  assign refill_full = (&{(! refill_slots_7_free),{(! refill_slots_6_free),{(! refill_slots_5_free),{(! refill_slots_4_free),{(! refill_slots_3_free),{(! refill_slots_2_free),{(! refill_slots_1_free),(! refill_slots_0_free)}}}}}}});
  always @(*) begin
    refill_push_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      refill_push_valid = 1'b1;
    end
    if(store_ctrl_startRefill) begin
      refill_push_valid = 1'b1;
    end
  end

  always @(*) begin
    refill_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(load_ctrl_startRefill) begin
      refill_push_payload_address = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
    end
    if(store_ctrl_startRefill) begin
      refill_push_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
    end
  end

  always @(*) begin
    refill_push_payload_way = 1'bx;
    refill_push_payload_way = load_ctrl_refillWay;
    if(store_ctrl_startRefill) begin
      refill_push_payload_way = store_ctrl_refillWay;
    end
  end

  always @(*) begin
    refill_push_payload_victim = 8'bxxxxxxxx;
    refill_push_payload_victim = ((load_ctrl_refillWayNeedWriteback && _zz_refill_push_payload_victim) ? writeback_free : 8'h0);
    if(store_ctrl_startRefill) begin
      refill_push_payload_victim = (((store_ctrl_replacedWayNeedWriteback && store_ctrl_askRefill) && _zz_refill_push_payload_victim_1) ? writeback_free : 8'h0);
    end
  end

  assign when_dcache2_l750 = refill_free[0];
  assign _zz_16 = refill_free[0];
  assign _zz_17 = refill_free[1];
  assign _zz_18 = refill_free[2];
  assign _zz_19 = refill_free[3];
  assign _zz_20 = refill_free[4];
  assign _zz_21 = refill_free[5];
  assign _zz_22 = refill_free[6];
  assign _zz_23 = refill_free[7];
  assign when_dcache2_l750_1 = refill_free[1];
  assign when_dcache2_l750_2 = refill_free[2];
  assign when_dcache2_l750_3 = refill_free[3];
  assign when_dcache2_l750_4 = refill_free[4];
  assign when_dcache2_l750_5 = refill_free[5];
  assign when_dcache2_l750_6 = refill_free[6];
  assign when_dcache2_l750_7 = refill_free[7];
  assign refill_read_arbiter_slotsWithId_0_0 = (((refill_slots_0_valid && (! refill_slots_0_cmdSent)) && (refill_slots_0_victim == 8'h0)) && (refill_slots_0_writebackHazards == 8'h0));
  assign refill_read_arbiter_slotsWithId_1_0 = (((refill_slots_1_valid && (! refill_slots_1_cmdSent)) && (refill_slots_1_victim == 8'h0)) && (refill_slots_1_writebackHazards == 8'h0));
  assign refill_read_arbiter_slotsWithId_2_0 = (((refill_slots_2_valid && (! refill_slots_2_cmdSent)) && (refill_slots_2_victim == 8'h0)) && (refill_slots_2_writebackHazards == 8'h0));
  assign refill_read_arbiter_slotsWithId_3_0 = (((refill_slots_3_valid && (! refill_slots_3_cmdSent)) && (refill_slots_3_victim == 8'h0)) && (refill_slots_3_writebackHazards == 8'h0));
  assign refill_read_arbiter_slotsWithId_4_0 = (((refill_slots_4_valid && (! refill_slots_4_cmdSent)) && (refill_slots_4_victim == 8'h0)) && (refill_slots_4_writebackHazards == 8'h0));
  assign refill_read_arbiter_slotsWithId_5_0 = (((refill_slots_5_valid && (! refill_slots_5_cmdSent)) && (refill_slots_5_victim == 8'h0)) && (refill_slots_5_writebackHazards == 8'h0));
  assign refill_read_arbiter_slotsWithId_6_0 = (((refill_slots_6_valid && (! refill_slots_6_cmdSent)) && (refill_slots_6_victim == 8'h0)) && (refill_slots_6_writebackHazards == 8'h0));
  assign refill_read_arbiter_slotsWithId_7_0 = (((refill_slots_7_valid && (! refill_slots_7_cmdSent)) && (refill_slots_7_victim == 8'h0)) && (refill_slots_7_writebackHazards == 8'h0));
  assign refill_read_arbiter_hits = {refill_read_arbiter_slotsWithId_7_0,{refill_read_arbiter_slotsWithId_6_0,{refill_read_arbiter_slotsWithId_5_0,{refill_read_arbiter_slotsWithId_4_0,{refill_read_arbiter_slotsWithId_3_0,{refill_read_arbiter_slotsWithId_2_0,{refill_read_arbiter_slotsWithId_1_0,refill_read_arbiter_slotsWithId_0_0}}}}}}};
  assign refill_read_arbiter_hit = (|refill_read_arbiter_hits);
  always @(*) begin
    refill_read_arbiter_oh = (refill_read_arbiter_hits & {(({_zz_refill_read_arbiter_oh,{_zz_refill_read_arbiter_oh_1,_zz_refill_read_arbiter_oh_2}} & refill_slots_7_priority) == 7'h0),{(({_zz_refill_read_arbiter_oh_9,_zz_refill_read_arbiter_oh_10} & refill_slots_6_priority) == 7'h0),{((_zz_refill_read_arbiter_oh_19 & refill_slots_5_priority) == 7'h0),{(_zz_refill_read_arbiter_oh_29 == _zz_refill_read_arbiter_oh_38),{_zz_refill_read_arbiter_oh_39,{_zz_refill_read_arbiter_oh_49,_zz_refill_read_arbiter_oh_60}}}}}});
    if(when_dcache2_l707) begin
      refill_read_arbiter_oh = refill_read_arbiter_lock;
    end
  end

  assign _zz_refill_read_arbiter_sel = refill_read_arbiter_oh[1];
  assign _zz_refill_read_arbiter_sel_1 = refill_read_arbiter_oh[2];
  assign _zz_refill_read_arbiter_sel_2 = refill_read_arbiter_oh[3];
  assign _zz_refill_read_arbiter_sel_3 = refill_read_arbiter_oh[4];
  assign _zz_refill_read_arbiter_sel_4 = refill_read_arbiter_oh[5];
  assign _zz_refill_read_arbiter_sel_5 = refill_read_arbiter_oh[6];
  assign _zz_refill_read_arbiter_sel_6 = refill_read_arbiter_oh[7];
  assign _zz_refill_read_arbiter_sel_7 = (((_zz_refill_read_arbiter_sel || _zz_refill_read_arbiter_sel_2) || _zz_refill_read_arbiter_sel_4) || _zz_refill_read_arbiter_sel_6);
  assign _zz_refill_read_arbiter_sel_8 = (((_zz_refill_read_arbiter_sel_1 || _zz_refill_read_arbiter_sel_2) || _zz_refill_read_arbiter_sel_5) || _zz_refill_read_arbiter_sel_6);
  assign _zz_refill_read_arbiter_sel_9 = (((_zz_refill_read_arbiter_sel_3 || _zz_refill_read_arbiter_sel_4) || _zz_refill_read_arbiter_sel_5) || _zz_refill_read_arbiter_sel_6);
  assign refill_read_arbiter_sel = {_zz_refill_read_arbiter_sel_9,{_zz_refill_read_arbiter_sel_8,_zz_refill_read_arbiter_sel_7}};
  assign when_dcache2_l707 = (|refill_read_arbiter_lock);
  assign refill_read_writebackHazard = (|refill_read_writebackHazards);
  assign io_mem_read_cmd_fire = (io_mem_read_cmd_valid && io_mem_read_cmd_ready);
  assign when_dcache2_l779 = (io_mem_read_cmd_fire || refill_read_writebackHazard);
  assign refill_read_cmdAddress = {_zz_refill_read_cmdAddress,5'h0};
  assign io_mem_read_cmd_valid = (refill_read_arbiter_hit && (! refill_read_writebackHazard));
  assign io_mem_read_cmd_payload_id = refill_read_arbiter_sel;
  assign io_mem_read_cmd_payload_address = refill_read_cmdAddress;
  assign when_dcache2_l791 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_dcache2_l791_1 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_dcache2_l791_2 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_dcache2_l791_3 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_dcache2_l791_4 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_dcache2_l791_5 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_dcache2_l791_6 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_dcache2_l791_7 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign refill_read_rspAddress = _zz_refill_read_rspAddress;
  assign refill_read_way = _zz_refill_read_way;
  assign refill_read_rspWithData = 1'b1;
  always @(*) begin
    refill_read_bankWriteNotif = 2'b00;
    refill_read_bankWriteNotif[0] = ((io_mem_read_rsp_valid && refill_read_rspWithData) && (refill_read_way == 1'b0));
    refill_read_bankWriteNotif[1] = ((io_mem_read_rsp_valid && refill_read_rspWithData) && (refill_read_way == 1'b1));
  end

  always @(*) begin
    banks_0_write_valid = refill_read_bankWriteNotif[0];
    if(store_ctrl_writeCache) begin
      if(when_dcache2_l1583) begin
        banks_0_write_valid = (1'b0 == store_ctrl_wayId);
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_address = {refill_read_rspAddress[8 : 5],refill_read_wordIndex};
    if(store_ctrl_writeCache) begin
      if(when_dcache2_l1583) begin
        banks_0_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 2];
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_data = io_mem_read_rsp_payload_data;
    if(store_ctrl_writeCache) begin
      if(when_dcache2_l1583) begin
        banks_0_write_payload_data[31 : 0] = store_pipeline_stages_2_CPU_WORD;
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_mask = 4'b1111;
    if(store_ctrl_writeCache) begin
      if(when_dcache2_l1583) begin
        banks_0_write_payload_mask = 4'b0000;
        if(_zz_when[0]) begin
          banks_0_write_payload_mask[3 : 0] = store_pipeline_stages_2_CPU_MASK;
        end
      end
    end
  end

  always @(*) begin
    banks_1_write_valid = refill_read_bankWriteNotif[1];
    if(store_ctrl_writeCache) begin
      if(when_dcache2_l1583_1) begin
        banks_1_write_valid = (1'b1 == store_ctrl_wayId);
      end
    end
  end

  always @(*) begin
    banks_1_write_payload_address = {refill_read_rspAddress[8 : 5],refill_read_wordIndex};
    if(store_ctrl_writeCache) begin
      if(when_dcache2_l1583_1) begin
        banks_1_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 2];
      end
    end
  end

  always @(*) begin
    banks_1_write_payload_data = io_mem_read_rsp_payload_data;
    if(store_ctrl_writeCache) begin
      if(when_dcache2_l1583_1) begin
        banks_1_write_payload_data[31 : 0] = store_pipeline_stages_2_CPU_WORD;
      end
    end
  end

  always @(*) begin
    banks_1_write_payload_mask = 4'b1111;
    if(store_ctrl_writeCache) begin
      if(when_dcache2_l1583_1) begin
        banks_1_write_payload_mask = 4'b0000;
        if(_zz_when_1[0]) begin
          banks_1_write_payload_mask[3 : 0] = store_pipeline_stages_2_CPU_MASK;
        end
      end
    end
  end

  assign when_dcache2_l821 = (io_mem_read_rsp_valid && io_mem_read_rsp_payload_error);
  always @(*) begin
    refill_read_fire = 1'b0;
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        refill_read_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    refill_read_reservation_take = 1'b0;
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        refill_read_reservation_take = 1'b1;
      end
    end
  end

  assign refill_read_faulty = (refill_read_hadError || io_mem_read_rsp_payload_error);
  always @(*) begin
    io_refillCompletions = 8'h0;
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        io_refillCompletions[io_mem_read_rsp_payload_id] = 1'b1;
      end
    end
  end

  assign io_mem_read_rsp_ready = 1'b1;
  assign when_dcache2_l834 = ((refill_read_wordIndex == 3'b111) || (! refill_read_rspWithData));
  always @(*) begin
    writeback_slots_0_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        3'b000 : begin
          writeback_slots_0_fire = 1'b1;
        end
        3'b001 : begin
        end
        3'b010 : begin
        end
        3'b011 : begin
        end
        3'b100 : begin
        end
        3'b101 : begin
        end
        3'b110 : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_0_free = (! writeback_slots_0_valid);
  always @(*) begin
    refill_read_writebackHazards[0] = (writeback_slots_0_valid && (writeback_slots_0_address[31 : 5] == refill_read_cmdAddress[31 : 5]));
    refill_read_writebackHazards[1] = (writeback_slots_1_valid && (writeback_slots_1_address[31 : 5] == refill_read_cmdAddress[31 : 5]));
    refill_read_writebackHazards[2] = (writeback_slots_2_valid && (writeback_slots_2_address[31 : 5] == refill_read_cmdAddress[31 : 5]));
    refill_read_writebackHazards[3] = (writeback_slots_3_valid && (writeback_slots_3_address[31 : 5] == refill_read_cmdAddress[31 : 5]));
    refill_read_writebackHazards[4] = (writeback_slots_4_valid && (writeback_slots_4_address[31 : 5] == refill_read_cmdAddress[31 : 5]));
    refill_read_writebackHazards[5] = (writeback_slots_5_valid && (writeback_slots_5_address[31 : 5] == refill_read_cmdAddress[31 : 5]));
    refill_read_writebackHazards[6] = (writeback_slots_6_valid && (writeback_slots_6_address[31 : 5] == refill_read_cmdAddress[31 : 5]));
    refill_read_writebackHazards[7] = (writeback_slots_7_valid && (writeback_slots_7_address[31 : 5] == refill_read_cmdAddress[31 : 5]));
  end

  always @(*) begin
    writeback_slots_1_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        3'b000 : begin
        end
        3'b001 : begin
          writeback_slots_1_fire = 1'b1;
        end
        3'b010 : begin
        end
        3'b011 : begin
        end
        3'b100 : begin
        end
        3'b101 : begin
        end
        3'b110 : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_1_free = (! writeback_slots_1_valid);
  always @(*) begin
    writeback_slots_2_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        3'b000 : begin
        end
        3'b001 : begin
        end
        3'b010 : begin
          writeback_slots_2_fire = 1'b1;
        end
        3'b011 : begin
        end
        3'b100 : begin
        end
        3'b101 : begin
        end
        3'b110 : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_2_free = (! writeback_slots_2_valid);
  always @(*) begin
    writeback_slots_3_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        3'b000 : begin
        end
        3'b001 : begin
        end
        3'b010 : begin
        end
        3'b011 : begin
          writeback_slots_3_fire = 1'b1;
        end
        3'b100 : begin
        end
        3'b101 : begin
        end
        3'b110 : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_3_free = (! writeback_slots_3_valid);
  always @(*) begin
    writeback_slots_4_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        3'b000 : begin
        end
        3'b001 : begin
        end
        3'b010 : begin
        end
        3'b011 : begin
        end
        3'b100 : begin
          writeback_slots_4_fire = 1'b1;
        end
        3'b101 : begin
        end
        3'b110 : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_4_free = (! writeback_slots_4_valid);
  always @(*) begin
    writeback_slots_5_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        3'b000 : begin
        end
        3'b001 : begin
        end
        3'b010 : begin
        end
        3'b011 : begin
        end
        3'b100 : begin
        end
        3'b101 : begin
          writeback_slots_5_fire = 1'b1;
        end
        3'b110 : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_5_free = (! writeback_slots_5_valid);
  always @(*) begin
    writeback_slots_6_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        3'b000 : begin
        end
        3'b001 : begin
        end
        3'b010 : begin
        end
        3'b011 : begin
        end
        3'b100 : begin
        end
        3'b101 : begin
        end
        3'b110 : begin
          writeback_slots_6_fire = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_6_free = (! writeback_slots_6_valid);
  always @(*) begin
    writeback_slots_7_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        3'b000 : begin
        end
        3'b001 : begin
        end
        3'b010 : begin
        end
        3'b011 : begin
        end
        3'b100 : begin
        end
        3'b101 : begin
        end
        3'b110 : begin
        end
        default : begin
          writeback_slots_7_fire = 1'b1;
        end
      endcase
    end
  end

  assign writeback_slots_7_free = (! writeback_slots_7_valid);
  assign io_writebackBusy = (|{writeback_slots_7_valid,{writeback_slots_6_valid,{writeback_slots_5_valid,{writeback_slots_4_valid,{writeback_slots_3_valid,{writeback_slots_2_valid,{writeback_slots_1_valid,writeback_slots_0_valid}}}}}}});
  assign _zz_writeback_free = {writeback_slots_7_free,{writeback_slots_6_free,{writeback_slots_5_free,{writeback_slots_4_free,{writeback_slots_3_free,{writeback_slots_2_free,{writeback_slots_1_free,writeback_slots_0_free}}}}}}};
  assign _zz_writeback_free_1 = (_zz_writeback_free & (~ _zz__zz_writeback_free_1));
  assign writeback_free = {_zz_writeback_free_1[7],{_zz_writeback_free_1[6],{_zz_writeback_free_1[5],{_zz_writeback_free_1[4],{_zz_writeback_free_1[3],{_zz_writeback_free_1[2],{_zz_writeback_free_1[1],writeback_slots_0_free}}}}}}};
  assign writeback_full = (&{(! writeback_slots_7_free),{(! writeback_slots_6_free),{(! writeback_slots_5_free),{(! writeback_slots_4_free),{(! writeback_slots_3_free),{(! writeback_slots_2_free),{(! writeback_slots_1_free),(! writeback_slots_0_free)}}}}}}});
  always @(*) begin
    writeback_push_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      writeback_push_valid = load_ctrl_refillWayNeedWriteback;
    end
    if(when_dcache2_l1552) begin
      writeback_push_valid = ((store_ctrl_replacedWayNeedWriteback && store_ctrl_startRefill) || store_ctrl_startFlush);
    end
  end

  always @(*) begin
    writeback_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(load_ctrl_startRefill) begin
      writeback_push_payload_address = ({5'd0,{_zz_writeback_push_payload_address,load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]}} <<< 3'd5);
    end
    if(when_dcache2_l1552) begin
      writeback_push_payload_address = ({5'd0,{_zz_writeback_push_payload_address_1,store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]}} <<< 3'd5);
    end
  end

  always @(*) begin
    writeback_push_payload_way = 1'bx;
    if(load_ctrl_startRefill) begin
      writeback_push_payload_way = load_ctrl_refillWay;
    end
    if(when_dcache2_l1552) begin
      writeback_push_payload_way = (store_pipeline_stages_2_FLUSH ? store_ctrl_needFlushSel : store_ctrl_refillWay);
    end
  end

  assign when_dcache2_l897 = writeback_free[0];
  assign _zz_24 = writeback_free[0];
  assign _zz_25 = writeback_free[1];
  assign _zz_26 = writeback_free[2];
  assign _zz_27 = writeback_free[3];
  assign _zz_28 = writeback_free[4];
  assign _zz_29 = writeback_free[5];
  assign _zz_30 = writeback_free[6];
  assign _zz_31 = writeback_free[7];
  assign when_dcache2_l897_1 = writeback_free[1];
  assign when_dcache2_l897_2 = writeback_free[2];
  assign when_dcache2_l897_3 = writeback_free[3];
  assign when_dcache2_l897_4 = writeback_free[4];
  assign when_dcache2_l897_5 = writeback_free[5];
  assign when_dcache2_l897_6 = writeback_free[6];
  assign when_dcache2_l897_7 = writeback_free[7];
  assign writeback_read_arbiter_slotsWithId_0_0 = (writeback_slots_0_valid && (! writeback_slots_0_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_1_0 = (writeback_slots_1_valid && (! writeback_slots_1_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_2_0 = (writeback_slots_2_valid && (! writeback_slots_2_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_3_0 = (writeback_slots_3_valid && (! writeback_slots_3_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_4_0 = (writeback_slots_4_valid && (! writeback_slots_4_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_5_0 = (writeback_slots_5_valid && (! writeback_slots_5_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_6_0 = (writeback_slots_6_valid && (! writeback_slots_6_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_7_0 = (writeback_slots_7_valid && (! writeback_slots_7_readCmdDone));
  assign writeback_read_arbiter_hits = {writeback_read_arbiter_slotsWithId_7_0,{writeback_read_arbiter_slotsWithId_6_0,{writeback_read_arbiter_slotsWithId_5_0,{writeback_read_arbiter_slotsWithId_4_0,{writeback_read_arbiter_slotsWithId_3_0,{writeback_read_arbiter_slotsWithId_2_0,{writeback_read_arbiter_slotsWithId_1_0,writeback_read_arbiter_slotsWithId_0_0}}}}}}};
  assign writeback_read_arbiter_hit = (|writeback_read_arbiter_hits);
  always @(*) begin
    writeback_read_arbiter_oh = (writeback_read_arbiter_hits & {(({_zz_writeback_read_arbiter_oh,{_zz_writeback_read_arbiter_oh_1,_zz_writeback_read_arbiter_oh_2}} & writeback_slots_7_priority) == 7'h0),{(({_zz_writeback_read_arbiter_oh_9,_zz_writeback_read_arbiter_oh_10} & writeback_slots_6_priority) == 7'h0),{((_zz_writeback_read_arbiter_oh_19 & writeback_slots_5_priority) == 7'h0),{(_zz_writeback_read_arbiter_oh_29 == _zz_writeback_read_arbiter_oh_38),{_zz_writeback_read_arbiter_oh_39,{_zz_writeback_read_arbiter_oh_49,_zz_writeback_read_arbiter_oh_60}}}}}});
    if(when_dcache2_l707_1) begin
      writeback_read_arbiter_oh = writeback_read_arbiter_lock;
    end
  end

  assign _zz_writeback_read_arbiter_sel = writeback_read_arbiter_oh[1];
  assign _zz_writeback_read_arbiter_sel_1 = writeback_read_arbiter_oh[2];
  assign _zz_writeback_read_arbiter_sel_2 = writeback_read_arbiter_oh[3];
  assign _zz_writeback_read_arbiter_sel_3 = writeback_read_arbiter_oh[4];
  assign _zz_writeback_read_arbiter_sel_4 = writeback_read_arbiter_oh[5];
  assign _zz_writeback_read_arbiter_sel_5 = writeback_read_arbiter_oh[6];
  assign _zz_writeback_read_arbiter_sel_6 = writeback_read_arbiter_oh[7];
  assign _zz_writeback_read_arbiter_sel_7 = (((_zz_writeback_read_arbiter_sel || _zz_writeback_read_arbiter_sel_2) || _zz_writeback_read_arbiter_sel_4) || _zz_writeback_read_arbiter_sel_6);
  assign _zz_writeback_read_arbiter_sel_8 = (((_zz_writeback_read_arbiter_sel_1 || _zz_writeback_read_arbiter_sel_2) || _zz_writeback_read_arbiter_sel_5) || _zz_writeback_read_arbiter_sel_6);
  assign _zz_writeback_read_arbiter_sel_9 = (((_zz_writeback_read_arbiter_sel_3 || _zz_writeback_read_arbiter_sel_4) || _zz_writeback_read_arbiter_sel_5) || _zz_writeback_read_arbiter_sel_6);
  assign writeback_read_arbiter_sel = {_zz_writeback_read_arbiter_sel_9,{_zz_writeback_read_arbiter_sel_8,_zz_writeback_read_arbiter_sel_7}};
  assign when_dcache2_l707_1 = (|writeback_read_arbiter_lock);
  assign writeback_read_address = _zz_writeback_read_address;
  assign writeback_read_way = _zz_writeback_read_way;
  assign writeback_read_slotRead_valid = writeback_read_arbiter_hit;
  assign writeback_read_slotRead_payload_id = writeback_read_arbiter_sel;
  assign writeback_read_slotRead_payload_wordIndex = writeback_read_wordIndex;
  assign writeback_read_slotRead_payload_way = writeback_read_way;
  assign writeback_read_slotRead_payload_last = (writeback_read_wordIndex == 3'b111);
  assign when_dcache2_l937 = (writeback_read_slotRead_valid && writeback_read_slotRead_payload_last);
  assign when_dcache2_l948 = (writeback_read_slotRead_valid && (writeback_read_way == 1'b0));
  assign when_dcache2_l948_1 = (writeback_read_slotRead_valid && (writeback_read_way == 1'b1));
  assign writeback_read_readedData = _zz_writeback_read_readedData;
  assign writeback_write_arbiter_slotsWithId_0_0 = ((writeback_slots_0_valid && writeback_slots_0_victimBufferReady) && (! writeback_slots_0_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_1_0 = ((writeback_slots_1_valid && writeback_slots_1_victimBufferReady) && (! writeback_slots_1_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_2_0 = ((writeback_slots_2_valid && writeback_slots_2_victimBufferReady) && (! writeback_slots_2_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_3_0 = ((writeback_slots_3_valid && writeback_slots_3_victimBufferReady) && (! writeback_slots_3_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_4_0 = ((writeback_slots_4_valid && writeback_slots_4_victimBufferReady) && (! writeback_slots_4_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_5_0 = ((writeback_slots_5_valid && writeback_slots_5_victimBufferReady) && (! writeback_slots_5_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_6_0 = ((writeback_slots_6_valid && writeback_slots_6_victimBufferReady) && (! writeback_slots_6_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_7_0 = ((writeback_slots_7_valid && writeback_slots_7_victimBufferReady) && (! writeback_slots_7_writeCmdDone));
  assign writeback_write_arbiter_hits = {writeback_write_arbiter_slotsWithId_7_0,{writeback_write_arbiter_slotsWithId_6_0,{writeback_write_arbiter_slotsWithId_5_0,{writeback_write_arbiter_slotsWithId_4_0,{writeback_write_arbiter_slotsWithId_3_0,{writeback_write_arbiter_slotsWithId_2_0,{writeback_write_arbiter_slotsWithId_1_0,writeback_write_arbiter_slotsWithId_0_0}}}}}}};
  assign writeback_write_arbiter_hit = (|writeback_write_arbiter_hits);
  always @(*) begin
    writeback_write_arbiter_oh = (writeback_write_arbiter_hits & {(({_zz_writeback_write_arbiter_oh,{_zz_writeback_write_arbiter_oh_1,_zz_writeback_write_arbiter_oh_2}} & writeback_slots_7_priority) == 7'h0),{(({_zz_writeback_write_arbiter_oh_9,_zz_writeback_write_arbiter_oh_10} & writeback_slots_6_priority) == 7'h0),{((_zz_writeback_write_arbiter_oh_19 & writeback_slots_5_priority) == 7'h0),{(_zz_writeback_write_arbiter_oh_29 == _zz_writeback_write_arbiter_oh_38),{_zz_writeback_write_arbiter_oh_39,{_zz_writeback_write_arbiter_oh_49,_zz_writeback_write_arbiter_oh_60}}}}}});
    if(when_dcache2_l707_2) begin
      writeback_write_arbiter_oh = writeback_write_arbiter_lock;
    end
  end

  assign _zz_writeback_write_arbiter_sel = writeback_write_arbiter_oh[1];
  assign _zz_writeback_write_arbiter_sel_1 = writeback_write_arbiter_oh[2];
  assign _zz_writeback_write_arbiter_sel_2 = writeback_write_arbiter_oh[3];
  assign _zz_writeback_write_arbiter_sel_3 = writeback_write_arbiter_oh[4];
  assign _zz_writeback_write_arbiter_sel_4 = writeback_write_arbiter_oh[5];
  assign _zz_writeback_write_arbiter_sel_5 = writeback_write_arbiter_oh[6];
  assign _zz_writeback_write_arbiter_sel_6 = writeback_write_arbiter_oh[7];
  assign _zz_writeback_write_arbiter_sel_7 = (((_zz_writeback_write_arbiter_sel || _zz_writeback_write_arbiter_sel_2) || _zz_writeback_write_arbiter_sel_4) || _zz_writeback_write_arbiter_sel_6);
  assign _zz_writeback_write_arbiter_sel_8 = (((_zz_writeback_write_arbiter_sel_1 || _zz_writeback_write_arbiter_sel_2) || _zz_writeback_write_arbiter_sel_5) || _zz_writeback_write_arbiter_sel_6);
  assign _zz_writeback_write_arbiter_sel_9 = (((_zz_writeback_write_arbiter_sel_3 || _zz_writeback_write_arbiter_sel_4) || _zz_writeback_write_arbiter_sel_5) || _zz_writeback_write_arbiter_sel_6);
  assign writeback_write_arbiter_sel = {_zz_writeback_write_arbiter_sel_9,{_zz_writeback_write_arbiter_sel_8,_zz_writeback_write_arbiter_sel_7}};
  assign when_dcache2_l707_2 = (|writeback_write_arbiter_lock);
  assign writeback_write_last = (writeback_write_wordIndex == 3'b111);
  assign writeback_write_bufferRead_valid = writeback_write_arbiter_hit;
  assign writeback_write_bufferRead_payload_id = writeback_write_arbiter_sel;
  assign writeback_write_bufferRead_payload_last = writeback_write_last;
  assign writeback_write_bufferRead_payload_address = _zz_writeback_write_bufferRead_payload_address;
  assign writeback_write_bufferRead_fire = (writeback_write_bufferRead_valid && writeback_write_bufferRead_ready);
  assign when_dcache2_l1020 = (writeback_write_bufferRead_fire && writeback_write_last);
  always @(*) begin
    writeback_write_bufferRead_ready = writeback_write_cmd_ready;
    if(when_Stream_l477) begin
      writeback_write_bufferRead_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! writeback_write_cmd_valid);
  assign writeback_write_cmd_valid = writeback_write_bufferRead_rValid;
  assign writeback_write_cmd_payload_id = writeback_write_bufferRead_rData_id;
  assign writeback_write_cmd_payload_address = writeback_write_bufferRead_rData_address;
  assign writeback_write_cmd_payload_last = writeback_write_bufferRead_rData_last;
  assign _zz_writeback_write_word = {writeback_write_bufferRead_payload_id,writeback_write_wordIndex};
  assign writeback_write_word = writeback_victimBuffer_spinal_port1;
  assign io_mem_write_cmd_valid = writeback_write_cmd_valid;
  assign writeback_write_cmd_ready = io_mem_write_cmd_ready;
  assign io_mem_write_cmd_payload_fragment_address = writeback_write_cmd_payload_address;
  assign io_mem_write_cmd_payload_fragment_data = writeback_write_word;
  assign io_mem_write_cmd_payload_fragment_id = writeback_write_cmd_payload_id;
  assign io_mem_write_cmd_payload_last = writeback_write_cmd_payload_last;
  assign _zz_load_pipeline_stages_0_throwRequest_dcache2_l1064 = io_load_cancels[0];
  assign load_pipeline_stages_0_throwRequest_dcache2_l1064 = _zz_load_pipeline_stages_0_throwRequest_dcache2_l1064;
  assign _zz_load_pipeline_stages_1_throwRequest_dcache2_l1064 = io_load_cancels[1];
  assign load_pipeline_stages_1_throwRequest_dcache2_l1064 = _zz_load_pipeline_stages_1_throwRequest_dcache2_l1064;
  assign load_pipeline_stages_2_throwRequest_dcache2_l1064 = io_load_cancels[2];
  assign load_pipeline_stages_1_WAYS_HAZARD_overloaded = (load_pipeline_stages_1_WAYS_HAZARD | ((waysWrite_addressLast == load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[8 : 5]) ? waysWrite_maskLast : 2'b00));
  assign io_load_cmd_ready = 1'b1;
  assign load_pipeline_stages_0_valid = io_load_cmd_valid;
  assign load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION = io_load_cmd_payload_virtual;
  assign load_pipeline_stages_0_REDO_ON_DATA_HAZARD = io_load_cmd_payload_redoOnDataHazard;
  assign load_pipeline_stages_0_TRANSACTION_ID = io_load_cmd_payload_id;
  assign load_pipeline_stages_0_WAYS_HAZARD = 2'b00;
  always @(*) begin
    load_pipeline_stages_0_BANK_BUSY[0] = banks_0_read_usedByWriteBack;
    load_pipeline_stages_0_BANK_BUSY[1] = banks_1_read_usedByWriteBack;
  end

  assign when_dcache2_l1108 = (! load_pipeline_stages_0_BANK_BUSY[0]);
  always @(*) begin
    load_pipeline_stages_0_BANK_BUSY_overloaded[0] = (load_pipeline_stages_0_BANK_BUSY[0] || (banks_0_write_valid && load_pipeline_stages_0_REDO_ON_DATA_HAZARD));
    load_pipeline_stages_0_BANK_BUSY_overloaded[1] = (load_pipeline_stages_0_BANK_BUSY[1] || (banks_1_write_valid && load_pipeline_stages_0_REDO_ON_DATA_HAZARD));
  end

  assign load_pipeline_stages_1_BANKS_WORDS_0 = banks_0_read_rsp;
  always @(*) begin
    load_pipeline_stages_1_BANK_BUSY_REMAPPED[0] = load_pipeline_stages_1_BANK_BUSY[1'b0];
    load_pipeline_stages_1_BANK_BUSY_REMAPPED[1] = load_pipeline_stages_1_BANK_BUSY[1'b1];
  end

  assign load_pipeline_stages_1_BANKS_MUXES_0 = load_pipeline_stages_1_BANKS_WORDS_0[31 : 0];
  assign when_dcache2_l1108_1 = (! load_pipeline_stages_0_BANK_BUSY[1]);
  assign load_pipeline_stages_1_BANKS_WORDS_1 = banks_1_read_rsp;
  assign load_pipeline_stages_1_BANKS_MUXES_1 = load_pipeline_stages_1_BANKS_WORDS_1[31 : 0];
  assign _zz_load_pipeline_stages_2_CPU_WORD = load_pipeline_stages_2_WAYS_HITS[1];
  assign load_pipeline_stages_2_CPU_WORD = ((load_pipeline_stages_2_WAYS_HITS[0] ? load_pipeline_stages_2_BANKS_MUXES_0 : 32'h0) | (_zz_load_pipeline_stages_2_CPU_WORD ? load_pipeline_stages_2_BANKS_MUXES_1 : 32'h0));
  assign load_pipeline_stages_0_ADDRESS_POST_TRANSLATION = io_load_translated_physical;
  assign load_pipeline_stages_0_ABORD = io_load_translated_abord;
  assign ways_0_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign ways_0_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[8 : 5];
  assign load_pipeline_stages_1_WAYS_TAGS_0_loaded = ways_0_loadRead_rsp_loaded;
  assign load_pipeline_stages_1_WAYS_TAGS_0_address = ways_0_loadRead_rsp_address;
  assign load_pipeline_stages_1_WAYS_TAGS_0_fault = ways_0_loadRead_rsp_fault;
  always @(*) begin
    load_pipeline_stages_1_WAYS_HITS[0] = (load_pipeline_stages_1_WAYS_TAGS_0_loaded && (load_pipeline_stages_1_WAYS_TAGS_0_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 9]));
    load_pipeline_stages_1_WAYS_HITS[1] = (load_pipeline_stages_1_WAYS_TAGS_1_loaded && (load_pipeline_stages_1_WAYS_TAGS_1_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 9]));
  end

  assign ways_1_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign ways_1_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[8 : 5];
  assign load_pipeline_stages_1_WAYS_TAGS_1_loaded = ways_1_loadRead_rsp_loaded;
  assign load_pipeline_stages_1_WAYS_TAGS_1_address = ways_1_loadRead_rsp_address;
  assign load_pipeline_stages_1_WAYS_TAGS_1_fault = ways_1_loadRead_rsp_fault;
  assign load_pipeline_stages_2_WAYS_HIT = (|load_pipeline_stages_2_WAYS_HITS);
  assign status_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign status_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[8 : 5];
  assign load_pipeline_stages_1_STATUS_0_dirty = status_loadRead_rsp_0_dirty;
  assign load_pipeline_stages_1_STATUS_1_dirty = status_loadRead_rsp_1_dirty;
  always @(*) begin
    _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = load_pipeline_stages_1_STATUS_0_dirty;
    if(when_dcache2_l659) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = status_writeLast_payload_data_0_dirty;
    end
    if(when_dcache2_l662) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = status_write_payload_data_0_dirty;
    end
  end

  always @(*) begin
    _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty = load_pipeline_stages_1_STATUS_1_dirty;
    if(when_dcache2_l659) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty = status_writeLast_payload_data_1_dirty;
    end
    if(when_dcache2_l662) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty = status_write_payload_data_1_dirty;
    end
  end

  assign when_dcache2_l659 = (status_writeLast_valid && (status_writeLast_payload_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[8 : 5]));
  assign when_dcache2_l662 = (status_write_valid && (status_write_payload_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[8 : 5]));
  assign load_pipeline_stages_1_STATUS_overloaded_0_dirty = _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  assign load_pipeline_stages_1_STATUS_overloaded_1_dirty = _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty;
  always @(*) begin
    load_pipeline_stages_1_REFILL_HITS_EARLY = {(refill_slots_7_valid && (refill_slots_7_address[31 : 5] == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5])),{(refill_slots_6_valid && (refill_slots_6_address[31 : 5] == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5])),{(refill_slots_5_valid && (_zz_load_pipeline_stages_1_REFILL_HITS_EARLY == _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_1)),{(refill_slots_4_valid && _zz_load_pipeline_stages_1_REFILL_HITS_EARLY_2),{_zz_load_pipeline_stages_1_REFILL_HITS_EARLY_3,{_zz_load_pipeline_stages_1_REFILL_HITS_EARLY_4,_zz_load_pipeline_stages_1_REFILL_HITS_EARLY_5}}}}}};
    if(load_refillCheckEarly_refillPushHit) begin
      if(_zz_16) begin
        load_pipeline_stages_1_REFILL_HITS_EARLY[0] = 1'b1;
      end
      if(_zz_17) begin
        load_pipeline_stages_1_REFILL_HITS_EARLY[1] = 1'b1;
      end
      if(_zz_18) begin
        load_pipeline_stages_1_REFILL_HITS_EARLY[2] = 1'b1;
      end
      if(_zz_19) begin
        load_pipeline_stages_1_REFILL_HITS_EARLY[3] = 1'b1;
      end
      if(_zz_20) begin
        load_pipeline_stages_1_REFILL_HITS_EARLY[4] = 1'b1;
      end
      if(_zz_21) begin
        load_pipeline_stages_1_REFILL_HITS_EARLY[5] = 1'b1;
      end
      if(_zz_22) begin
        load_pipeline_stages_1_REFILL_HITS_EARLY[6] = 1'b1;
      end
      if(_zz_23) begin
        load_pipeline_stages_1_REFILL_HITS_EARLY[7] = 1'b1;
      end
    end
  end

  assign load_refillCheckEarly_refillPushHit = (refill_push_valid && (refill_push_payload_address[31 : 5] == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]));
  assign load_pipeline_stages_2_REFILL_HITS = (load_pipeline_stages_2_REFILL_HITS_EARLY & {refill_slots_7_valid,{refill_slots_6_valid,{refill_slots_5_valid,{refill_slots_4_valid,{refill_slots_3_valid,{refill_slots_2_valid,{refill_slots_1_valid,refill_slots_0_valid}}}}}}});
  always @(*) begin
    load_ctrl_reservation_take = 1'b0;
    if(load_ctrl_startRefill) begin
      load_ctrl_reservation_take = 1'b1;
    end
  end

  assign load_ctrl_refillWay = wayRandom_value;
  assign _zz_refill_push_payload_victim = _zz__zz_refill_push_payload_victim;
  assign load_ctrl_refillWayNeedWriteback = (_zz_load_ctrl_refillWayNeedWriteback && _zz_refill_push_payload_victim);
  assign load_ctrl_refillHit = (|load_pipeline_stages_2_REFILL_HITS);
  assign load_ctrl_refillLoaded = (|({refill_slots_7_loaded,{refill_slots_6_loaded,{refill_slots_5_loaded,{refill_slots_4_loaded,{refill_slots_3_loaded,{refill_slots_2_loaded,{refill_slots_1_loaded,refill_slots_0_loaded}}}}}}} & load_pipeline_stages_2_REFILL_HITS));
  assign load_ctrl_lineBusy = ((|{(refill_slots_7_valid && (_zz_load_ctrl_lineBusy == _zz_load_ctrl_lineBusy_1)),{(refill_slots_6_valid && _zz_load_ctrl_lineBusy_2),{_zz_load_ctrl_lineBusy_3,{_zz_load_ctrl_lineBusy_6,_zz_load_ctrl_lineBusy_8}}}}) || (|{(writeback_slots_7_valid && (_zz_load_ctrl_lineBusy_16 == _zz_load_ctrl_lineBusy_17)),{(writeback_slots_6_valid && _zz_load_ctrl_lineBusy_18),{_zz_load_ctrl_lineBusy_19,{_zz_load_ctrl_lineBusy_22,_zz_load_ctrl_lineBusy_24}}}}));
  assign load_ctrl_bankBusy = ((load_pipeline_stages_2_BANK_BUSY_REMAPPED & load_pipeline_stages_2_WAYS_HITS) != 2'b00);
  assign load_ctrl_waysHitHazard = (|(load_pipeline_stages_2_WAYS_HITS & load_pipeline_stages_2_WAYS_HAZARD_resulting));
  always @(*) begin
    load_pipeline_stages_2_REDO = ((((! load_pipeline_stages_2_WAYS_HIT) || load_ctrl_waysHitHazard) || load_ctrl_bankBusy) || load_ctrl_refillHit);
    if(load_pipeline_stages_2_ABORD) begin
      load_pipeline_stages_2_REDO = 1'b0;
    end
  end

  always @(*) begin
    load_pipeline_stages_2_MISS = (((! load_pipeline_stages_2_WAYS_HIT) && (! load_ctrl_waysHitHazard)) && (! load_ctrl_refillHit));
    if(load_pipeline_stages_2_ABORD) begin
      load_pipeline_stages_2_MISS = 1'b0;
    end
  end

  assign load_pipeline_stages_2_FAULT = (|(load_pipeline_stages_2_WAYS_HITS & {load_pipeline_stages_2_WAYS_TAGS_1_fault,load_pipeline_stages_2_WAYS_TAGS_0_fault}));
  assign load_ctrl_canRefill = (((((! refill_full) && (! load_ctrl_lineBusy)) && load_ctrl_reservation_win) && (! (load_ctrl_refillWayNeedWriteback && writeback_full))) && (! load_pipeline_stages_2_WAYS_HAZARD_resulting[load_ctrl_refillWay]));
  assign load_ctrl_askRefill = ((load_pipeline_stages_2_MISS && load_ctrl_canRefill) && (! load_ctrl_refillHit));
  assign load_ctrl_startRefill = (load_pipeline_stages_2_valid && load_ctrl_askRefill);
  assign load_ctrl_wayId = _zz_load_pipeline_stages_2_CPU_WORD;
  assign _zz_34 = ({1'd0,1'b1} <<< load_ctrl_refillWay);
  assign load_pipeline_stages_2_REFILL_SLOT_FULL = ((load_pipeline_stages_2_MISS && (! load_ctrl_refillHit)) && refill_full);
  assign load_pipeline_stages_2_REFILL_SLOT = (((! load_ctrl_refillLoaded) ? load_pipeline_stages_2_REFILL_HITS : 8'h0) | (load_ctrl_askRefill ? refill_free : 8'h0));
  assign io_load_rsp_valid = load_pipeline_stages_2_valid;
  assign io_load_rsp_payload_data = load_pipeline_stages_2_CPU_WORD;
  assign io_load_rsp_payload_fault = load_pipeline_stages_2_FAULT;
  assign io_load_rsp_payload_redo = load_pipeline_stages_2_REDO;
  assign io_load_rsp_payload_id = load_pipeline_stages_2_TRANSACTION_ID;
  assign io_load_rsp_payload_refillSlotAny = load_pipeline_stages_2_REFILL_SLOT_FULL;
  assign io_load_rsp_payload_refillSlot = load_pipeline_stages_2_REFILL_SLOT;
  assign load_pipeline_stages_2_isThrown = load_pipeline_stages_2_throwRequest_dcache2_l1064;
  assign load_pipeline_stages_1_isThrown = load_pipeline_stages_1_throwRequest_dcache2_l1064;
  assign load_pipeline_stages_0_isThrown = load_pipeline_stages_0_throwRequest_dcache2_l1064;
  always @(*) begin
    _zz_load_pipeline_stages_1_valid = load_pipeline_stages_0_valid;
    if(when_Pipeline_l276) begin
      _zz_load_pipeline_stages_1_valid = 1'b0;
    end
  end

  assign load_pipeline_stages_0_ready = 1'b1;
  assign when_Pipeline_l276 = (|_zz_load_pipeline_stages_0_throwRequest_dcache2_l1064);
  always @(*) begin
    _zz_load_pipeline_stages_2_valid = load_pipeline_stages_1_valid;
    if(when_Pipeline_l276_1) begin
      _zz_load_pipeline_stages_2_valid = 1'b0;
    end
  end

  assign load_pipeline_stages_1_ready = 1'b1;
  assign when_Pipeline_l276_1 = (|_zz_load_pipeline_stages_1_throwRequest_dcache2_l1064);
  assign load_pipeline_stages_2_WAYS_HAZARD_resulting = load_pipeline_stages_2_WAYS_HAZARD;
  assign store_pipeline_discardAll = 1'b0;
  assign store_pipeline_stages_0_throwRequest_dcache2_l1357 = store_pipeline_discardAll;
  assign store_pipeline_stages_1_throwRequest_dcache2_l1357 = store_pipeline_discardAll;
  assign store_pipeline_stages_2_throwRequest_dcache2_l1357 = store_pipeline_discardAll;
  assign store_pipeline_stages_1_WAYS_HAZARD_overloaded = (store_pipeline_stages_1_WAYS_HAZARD | ((waysWrite_addressLast == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[8 : 5]) ? waysWrite_maskLast : 2'b00));
  assign store_pipeline_stages_2_WAYS_HAZARD_overloaded = (store_pipeline_stages_2_WAYS_HAZARD | ((waysWrite_addressLast == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5]) ? waysWrite_maskLast : 2'b00));
  assign store_pipeline_stages_0_valid = io_store_cmd_valid;
  assign store_pipeline_stages_0_ADDRESS_POST_TRANSLATION = io_store_cmd_payload_address;
  assign store_pipeline_stages_0_CPU_WORD = io_store_cmd_payload_data;
  assign store_pipeline_stages_0_CPU_MASK = io_store_cmd_payload_mask;
  assign store_pipeline_stages_0_IO = (io_store_cmd_payload_io && (! io_store_cmd_payload_flush));
  assign store_pipeline_stages_0_FLUSH = io_store_cmd_payload_flush;
  assign store_pipeline_stages_0_FLUSH_FREE = io_store_cmd_payload_flushFree;
  assign store_pipeline_stages_0_PREFETCH = io_store_cmd_payload_prefetch;
  assign store_pipeline_stages_0_TRANSACTION_ID = io_store_cmd_payload_id;
  assign store_pipeline_stages_0_WAYS_HAZARD = 2'b00;
  assign io_store_cmd_ready = 1'b1;
  assign ways_0_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign ways_0_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[8 : 5];
  assign store_pipeline_stages_1_WAYS_TAGS_0_loaded = ways_0_storeRead_rsp_loaded;
  assign store_pipeline_stages_1_WAYS_TAGS_0_address = ways_0_storeRead_rsp_address;
  assign store_pipeline_stages_1_WAYS_TAGS_0_fault = ways_0_storeRead_rsp_fault;
  always @(*) begin
    store_pipeline_stages_1_WAYS_HITS[0] = (store_pipeline_stages_1_WAYS_TAGS_0_loaded && (store_pipeline_stages_1_WAYS_TAGS_0_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 9]));
    store_pipeline_stages_1_WAYS_HITS[1] = (store_pipeline_stages_1_WAYS_TAGS_1_loaded && (store_pipeline_stages_1_WAYS_TAGS_1_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 9]));
  end

  assign _zz_35 = store_pipeline_stages_1_WAYS_HITS[0];
  assign ways_1_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign ways_1_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[8 : 5];
  assign store_pipeline_stages_1_WAYS_TAGS_1_loaded = ways_1_storeRead_rsp_loaded;
  assign store_pipeline_stages_1_WAYS_TAGS_1_address = ways_1_storeRead_rsp_address;
  assign store_pipeline_stages_1_WAYS_TAGS_1_fault = ways_1_storeRead_rsp_fault;
  assign _zz_36 = store_pipeline_stages_1_WAYS_HITS[1];
  assign store_pipeline_stages_1_WAYS_HIT = (|store_pipeline_stages_1_WAYS_HITS);
  assign _zz_37 = store_pipeline_stages_1_WAYS_HIT;
  assign _zz_38 = store_pipeline_stages_1_WAYS_HITS;
  assign status_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign status_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[8 : 5];
  assign store_pipeline_stages_1_STATUS_0_dirty = status_storeRead_rsp_0_dirty;
  assign store_pipeline_stages_1_STATUS_1_dirty = status_storeRead_rsp_1_dirty;
  always @(*) begin
    _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = store_pipeline_stages_1_STATUS_0_dirty;
    if(when_dcache2_l659_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = status_writeLast_payload_data_0_dirty;
    end
    if(when_dcache2_l662_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = status_write_payload_data_0_dirty;
    end
  end

  always @(*) begin
    _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty = store_pipeline_stages_1_STATUS_1_dirty;
    if(when_dcache2_l659_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty = status_writeLast_payload_data_1_dirty;
    end
    if(when_dcache2_l662_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty = status_write_payload_data_1_dirty;
    end
  end

  assign when_dcache2_l659_1 = (status_writeLast_valid && (status_writeLast_payload_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[8 : 5]));
  assign when_dcache2_l662_1 = (status_write_valid && (status_write_payload_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[8 : 5]));
  assign store_pipeline_stages_1_STATUS_overloaded_0_dirty = _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  assign store_pipeline_stages_1_STATUS_overloaded_1_dirty = _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty;
  always @(*) begin
    store_pipeline_stages_1_REFILL_HITS_EARLY = {(refill_slots_7_valid && (refill_slots_7_address[31 : 5] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5])),{(refill_slots_6_valid && (refill_slots_6_address[31 : 5] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5])),{(refill_slots_5_valid && (_zz_store_pipeline_stages_1_REFILL_HITS_EARLY == _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_1)),{(refill_slots_4_valid && _zz_store_pipeline_stages_1_REFILL_HITS_EARLY_2),{_zz_store_pipeline_stages_1_REFILL_HITS_EARLY_3,{_zz_store_pipeline_stages_1_REFILL_HITS_EARLY_4,_zz_store_pipeline_stages_1_REFILL_HITS_EARLY_5}}}}}};
    if(store_refillCheckEarly_refillPushHit) begin
      if(_zz_16) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[0] = 1'b1;
      end
      if(_zz_17) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[1] = 1'b1;
      end
      if(_zz_18) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[2] = 1'b1;
      end
      if(_zz_19) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[3] = 1'b1;
      end
      if(_zz_20) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[4] = 1'b1;
      end
      if(_zz_21) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[5] = 1'b1;
      end
      if(_zz_22) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[6] = 1'b1;
      end
      if(_zz_23) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[7] = 1'b1;
      end
    end
  end

  assign store_refillCheckEarly_refillPushHit = (refill_push_valid && (refill_push_payload_address[31 : 5] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 5]));
  assign store_pipeline_stages_2_REFILL_HITS = (store_pipeline_stages_2_REFILL_HITS_EARLY & {refill_slots_7_valid,{refill_slots_6_valid,{refill_slots_5_valid,{refill_slots_4_valid,{refill_slots_3_valid,{refill_slots_2_valid,{refill_slots_1_valid,refill_slots_0_valid}}}}}}});
  assign store_ctrl_generationOk = 1'b1;
  always @(*) begin
    store_ctrl_reservation_take = 1'b0;
    if(when_dcache2_l1542) begin
      store_ctrl_reservation_take = 1'b1;
    end
  end

  assign store_ctrl_replacedWay = wayRandom_value;
  assign store_ctrl_replacedWayNeedWriteback = (_zz_store_ctrl_replacedWayNeedWriteback && _zz_store_ctrl_replacedWayNeedWriteback_1);
  assign store_ctrl_refillHit = (|(store_pipeline_stages_2_REFILL_HITS & {refill_slots_7_valid,{refill_slots_6_valid,{refill_slots_5_valid,{refill_slots_4_valid,{refill_slots_3_valid,{refill_slots_2_valid,{refill_slots_1_valid,refill_slots_0_valid}}}}}}}));
  assign store_ctrl_lineBusy = ((|{(refill_slots_7_valid && (_zz_store_ctrl_lineBusy == _zz_store_ctrl_lineBusy_1)),{(refill_slots_6_valid && _zz_store_ctrl_lineBusy_2),{_zz_store_ctrl_lineBusy_3,{_zz_store_ctrl_lineBusy_6,_zz_store_ctrl_lineBusy_8}}}}) || (|{(writeback_slots_7_valid && (_zz_store_ctrl_lineBusy_16 == _zz_store_ctrl_lineBusy_17)),{(writeback_slots_6_valid && _zz_store_ctrl_lineBusy_18),{_zz_store_ctrl_lineBusy_19,{_zz_store_ctrl_lineBusy_22,_zz_store_ctrl_lineBusy_24}}}}));
  assign store_ctrl_waysHitHazard = (|(store_pipeline_stages_2_WAYS_HITS & store_pipeline_stages_2_WAYS_HAZARD_resulting));
  assign store_ctrl_wasClean = (! (|({store_pipeline_stages_2_STATUS_1_dirty,store_pipeline_stages_2_STATUS_0_dirty} & store_pipeline_stages_2_WAYS_HITS)));
  assign store_ctrl_bankBusy = (((! store_pipeline_stages_2_FLUSH) && (! store_pipeline_stages_2_PREFETCH)) && (|(store_pipeline_stages_2_WAYS_HITS & refill_read_bankWriteNotif)));
  assign store_ctrl_hitFault = (|(store_pipeline_stages_2_WAYS_HITS & {store_pipeline_stages_2_WAYS_TAGS_1_fault,store_pipeline_stages_2_WAYS_TAGS_0_fault}));
  assign store_ctrl_refillWay = store_ctrl_replacedWay;
  always @(*) begin
    store_pipeline_stages_2_REDO = (((((store_pipeline_stages_2_MISS || store_ctrl_waysHitHazard) || store_ctrl_bankBusy) || store_ctrl_refillHit) || (! store_ctrl_generationOk)) || (store_ctrl_wasClean && (! store_ctrl_reservation_win)));
    if(store_pipeline_stages_2_FLUSH) begin
      store_pipeline_stages_2_REDO = (store_ctrl_needFlush || (|store_pipeline_stages_2_WAYS_HAZARD_resulting));
    end
    if(store_pipeline_stages_2_IO) begin
      store_pipeline_stages_2_REDO = 1'b0;
    end
  end

  always @(*) begin
    store_pipeline_stages_2_MISS = (((! store_pipeline_stages_2_WAYS_HIT) && (! store_ctrl_waysHitHazard)) && (! store_ctrl_refillHit));
    if(store_pipeline_stages_2_IO) begin
      store_pipeline_stages_2_MISS = 1'b0;
    end
  end

  assign store_ctrl_canRefill = (((((! refill_full) && (! store_ctrl_lineBusy)) && (! load_ctrl_startRefill)) && store_ctrl_reservation_win) && (! store_pipeline_stages_2_WAYS_HAZARD_resulting[store_ctrl_refillWay]));
  assign store_ctrl_askRefill = (((store_pipeline_stages_2_MISS && store_ctrl_canRefill) && (! store_ctrl_refillHit)) && (! (store_ctrl_replacedWayNeedWriteback && writeback_full)));
  always @(*) begin
    store_ctrl_startRefill = ((store_pipeline_stages_2_valid && store_ctrl_generationOk) && store_ctrl_askRefill);
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_startRefill = 1'b0;
    end
  end

  assign store_pipeline_stages_2_REFILL_SLOT_FULL = ((store_pipeline_stages_2_MISS && (! store_ctrl_refillHit)) && refill_full);
  assign store_pipeline_stages_2_REFILL_SLOT = (store_ctrl_askRefill ? refill_free : 8'h0);
  always @(*) begin
    store_ctrl_writeCache = (((store_pipeline_stages_2_valid && store_ctrl_generationOk) && (! store_pipeline_stages_2_REDO)) && (! store_pipeline_stages_2_PREFETCH));
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_writeCache = 1'b0;
    end
    if(store_pipeline_stages_2_IO) begin
      store_ctrl_writeCache = 1'b0;
    end
  end

  always @(*) begin
    store_ctrl_setDirty = (store_ctrl_writeCache && store_ctrl_wasClean);
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_setDirty = 1'b0;
    end
    if(store_pipeline_stages_2_IO) begin
      store_ctrl_setDirty = 1'b0;
    end
  end

  assign _zz_store_ctrl_wayId = store_pipeline_stages_2_WAYS_HITS[1];
  assign store_ctrl_wayId = _zz_store_ctrl_wayId;
  assign store_ctrl_needFlushs = ({store_pipeline_stages_2_WAYS_TAGS_1_loaded,store_pipeline_stages_2_WAYS_TAGS_0_loaded} & {store_pipeline_stages_2_STATUS_1_dirty,store_pipeline_stages_2_STATUS_0_dirty});
  assign _zz_store_ctrl_needFlushs_bools_0 = store_ctrl_needFlushs;
  assign store_ctrl_needFlushs_bools_0 = _zz_store_ctrl_needFlushs_bools_0[0];
  assign store_ctrl_needFlushs_bools_1 = _zz_store_ctrl_needFlushs_bools_0[1];
  always @(*) begin
    _zz_store_ctrl_needFlushOh[0] = (store_ctrl_needFlushs_bools_0 && (! 1'b0));
    _zz_store_ctrl_needFlushOh[1] = (store_ctrl_needFlushs_bools_1 && (! store_ctrl_needFlushs_bools_0));
  end

  assign store_ctrl_needFlushOh = _zz_store_ctrl_needFlushOh;
  assign _zz_store_ctrl_needFlushSel = store_ctrl_needFlushOh[1];
  assign store_ctrl_needFlushSel = _zz_store_ctrl_needFlushSel;
  assign store_ctrl_needFlush = (|store_ctrl_needFlushs);
  assign store_ctrl_canFlush = (((store_ctrl_reservation_win && (! writeback_full)) && (! (|{refill_slots_7_valid,{refill_slots_6_valid,{refill_slots_5_valid,{refill_slots_4_valid,{refill_slots_3_valid,{refill_slots_2_valid,{refill_slots_1_valid,refill_slots_0_valid}}}}}}}))) && (! (|store_pipeline_stages_2_WAYS_HAZARD_resulting)));
  assign store_ctrl_startFlush = ((((store_pipeline_stages_2_valid && store_pipeline_stages_2_FLUSH) && store_ctrl_generationOk) && store_ctrl_needFlush) && store_ctrl_canFlush);
  assign when_dcache2_l1542 = ((store_ctrl_startRefill || store_ctrl_setDirty) || store_ctrl_startFlush);
  assign when_dcache2_l1552 = (store_ctrl_startRefill || store_ctrl_startFlush);
  assign when_dcache2_l1583 = store_pipeline_stages_2_WAYS_HITS[0];
  assign when_dcache2_l1583_1 = store_pipeline_stages_2_WAYS_HITS[1];
  assign _zz_40 = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_41 = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[8 : 5];
  assign _zz_42 = store_pipeline_stages_2_WAYS_HIT;
  assign _zz_43 = store_pipeline_stages_2_MISS;
  assign _zz_44 = store_pipeline_stages_2_REDO;
  assign _zz_45 = store_pipeline_stages_2_IO;
  assign _zz_46 = store_pipeline_stages_2_FLUSH;
  assign _zz_47 = store_pipeline_stages_2_PREFETCH;
  assign io_store_rsp_valid = store_pipeline_stages_2_valid;
  assign io_store_rsp_payload_fault = 1'b0;
  assign io_store_rsp_payload_redo = store_pipeline_stages_2_REDO;
  assign io_store_rsp_payload_id = store_pipeline_stages_2_TRANSACTION_ID;
  assign io_store_rsp_payload_refillSlotAny = store_pipeline_stages_2_REFILL_SLOT_FULL;
  assign io_store_rsp_payload_refillSlot = store_pipeline_stages_2_REFILL_SLOT;
  assign io_store_rsp_payload_flush = store_pipeline_stages_2_FLUSH;
  assign io_store_rsp_payload_prefetch = store_pipeline_stages_2_PREFETCH;
  assign io_store_rsp_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  assign io_store_rsp_payload_io = store_pipeline_stages_2_IO;
  assign store_pipeline_stages_2_isThrown = store_pipeline_stages_2_throwRequest_dcache2_l1357;
  assign store_pipeline_stages_1_isThrown = store_pipeline_stages_1_throwRequest_dcache2_l1357;
  assign store_pipeline_stages_0_isThrown = store_pipeline_stages_0_throwRequest_dcache2_l1357;
  always @(*) begin
    _zz_store_pipeline_stages_1_valid = store_pipeline_stages_0_valid;
    if(when_Pipeline_l276_2) begin
      _zz_store_pipeline_stages_1_valid = 1'b0;
    end
  end

  assign when_Pipeline_l276_2 = (|store_pipeline_discardAll);
  always @(*) begin
    _zz_store_pipeline_stages_2_valid = store_pipeline_stages_1_valid;
    if(when_Pipeline_l276_3) begin
      _zz_store_pipeline_stages_2_valid = 1'b0;
    end
  end

  assign store_pipeline_stages_1_ready = 1'b1;
  assign when_Pipeline_l276_3 = (|store_pipeline_discardAll);
  assign store_pipeline_stages_2_WAYS_HAZARD_resulting = store_pipeline_stages_2_WAYS_HAZARD_overloaded;
  assign io_refillEvent = refill_push_valid;
  assign io_writebackEvent = writeback_push_valid;
  assign invalidate_reservation_win = (! 1'b0);
  assign refill_read_reservation_win = (! 1'b0);
  assign load_ctrl_reservation_win = (! (|{refill_read_reservation_take,invalidate_reservation_take}));
  assign store_ctrl_reservation_win = (! (|{load_ctrl_reservation_take,{refill_read_reservation_take,invalidate_reservation_take}}));
  always @(posedge clk) begin
    waysWrite_maskLast <= waysWrite_mask;
    waysWrite_addressLast <= waysWrite_address;
    status_writeLast_payload_address <= status_write_payload_address;
    status_writeLast_payload_data_0_dirty <= status_write_payload_data_0_dirty;
    status_writeLast_payload_data_1_dirty <= status_write_payload_data_1_dirty;
    refill_slots_0_loadedCounter <= (refill_slots_0_loadedCounter + (refill_slots_0_loaded && (! refill_slots_0_loadedDone)));
    refill_slots_1_loadedCounter <= (refill_slots_1_loadedCounter + (refill_slots_1_loaded && (! refill_slots_1_loadedDone)));
    refill_slots_2_loadedCounter <= (refill_slots_2_loadedCounter + (refill_slots_2_loaded && (! refill_slots_2_loadedDone)));
    refill_slots_3_loadedCounter <= (refill_slots_3_loadedCounter + (refill_slots_3_loaded && (! refill_slots_3_loadedDone)));
    refill_slots_4_loadedCounter <= (refill_slots_4_loadedCounter + (refill_slots_4_loaded && (! refill_slots_4_loadedDone)));
    refill_slots_5_loadedCounter <= (refill_slots_5_loadedCounter + (refill_slots_5_loaded && (! refill_slots_5_loadedDone)));
    refill_slots_6_loadedCounter <= (refill_slots_6_loadedCounter + (refill_slots_6_loaded && (! refill_slots_6_loadedDone)));
    refill_slots_7_loadedCounter <= (refill_slots_7_loadedCounter + (refill_slots_7_loaded && (! refill_slots_7_loadedDone)));
    if(refill_push_valid) begin
      if(when_dcache2_l750) begin
        refill_slots_0_address <= refill_push_payload_address;
        refill_slots_0_way <= refill_push_payload_way;
        refill_slots_0_cmdSent <= 1'b0;
        refill_slots_0_priority <= 7'h7f;
        refill_slots_0_loaded <= 1'b0;
        refill_slots_0_loadedCounter <= 1'b0;
        refill_slots_0_victim <= refill_push_payload_victim;
        refill_slots_0_writebackHazards <= 8'h0;
      end else begin
        if(_zz_17) begin
          refill_slots_0_priority[0] <= 1'b0;
        end
        if(_zz_18) begin
          refill_slots_0_priority[1] <= 1'b0;
        end
        if(_zz_19) begin
          refill_slots_0_priority[2] <= 1'b0;
        end
        if(_zz_20) begin
          refill_slots_0_priority[3] <= 1'b0;
        end
        if(_zz_21) begin
          refill_slots_0_priority[4] <= 1'b0;
        end
        if(_zz_22) begin
          refill_slots_0_priority[5] <= 1'b0;
        end
        if(_zz_23) begin
          refill_slots_0_priority[6] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_dcache2_l750_1) begin
        refill_slots_1_address <= refill_push_payload_address;
        refill_slots_1_way <= refill_push_payload_way;
        refill_slots_1_cmdSent <= 1'b0;
        refill_slots_1_priority <= 7'h7f;
        refill_slots_1_loaded <= 1'b0;
        refill_slots_1_loadedCounter <= 1'b0;
        refill_slots_1_victim <= refill_push_payload_victim;
        refill_slots_1_writebackHazards <= 8'h0;
      end else begin
        if(_zz_16) begin
          refill_slots_1_priority[0] <= 1'b0;
        end
        if(_zz_18) begin
          refill_slots_1_priority[1] <= 1'b0;
        end
        if(_zz_19) begin
          refill_slots_1_priority[2] <= 1'b0;
        end
        if(_zz_20) begin
          refill_slots_1_priority[3] <= 1'b0;
        end
        if(_zz_21) begin
          refill_slots_1_priority[4] <= 1'b0;
        end
        if(_zz_22) begin
          refill_slots_1_priority[5] <= 1'b0;
        end
        if(_zz_23) begin
          refill_slots_1_priority[6] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_dcache2_l750_2) begin
        refill_slots_2_address <= refill_push_payload_address;
        refill_slots_2_way <= refill_push_payload_way;
        refill_slots_2_cmdSent <= 1'b0;
        refill_slots_2_priority <= 7'h7f;
        refill_slots_2_loaded <= 1'b0;
        refill_slots_2_loadedCounter <= 1'b0;
        refill_slots_2_victim <= refill_push_payload_victim;
        refill_slots_2_writebackHazards <= 8'h0;
      end else begin
        if(_zz_16) begin
          refill_slots_2_priority[0] <= 1'b0;
        end
        if(_zz_17) begin
          refill_slots_2_priority[1] <= 1'b0;
        end
        if(_zz_19) begin
          refill_slots_2_priority[2] <= 1'b0;
        end
        if(_zz_20) begin
          refill_slots_2_priority[3] <= 1'b0;
        end
        if(_zz_21) begin
          refill_slots_2_priority[4] <= 1'b0;
        end
        if(_zz_22) begin
          refill_slots_2_priority[5] <= 1'b0;
        end
        if(_zz_23) begin
          refill_slots_2_priority[6] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_dcache2_l750_3) begin
        refill_slots_3_address <= refill_push_payload_address;
        refill_slots_3_way <= refill_push_payload_way;
        refill_slots_3_cmdSent <= 1'b0;
        refill_slots_3_priority <= 7'h7f;
        refill_slots_3_loaded <= 1'b0;
        refill_slots_3_loadedCounter <= 1'b0;
        refill_slots_3_victim <= refill_push_payload_victim;
        refill_slots_3_writebackHazards <= 8'h0;
      end else begin
        if(_zz_16) begin
          refill_slots_3_priority[0] <= 1'b0;
        end
        if(_zz_17) begin
          refill_slots_3_priority[1] <= 1'b0;
        end
        if(_zz_18) begin
          refill_slots_3_priority[2] <= 1'b0;
        end
        if(_zz_20) begin
          refill_slots_3_priority[3] <= 1'b0;
        end
        if(_zz_21) begin
          refill_slots_3_priority[4] <= 1'b0;
        end
        if(_zz_22) begin
          refill_slots_3_priority[5] <= 1'b0;
        end
        if(_zz_23) begin
          refill_slots_3_priority[6] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_dcache2_l750_4) begin
        refill_slots_4_address <= refill_push_payload_address;
        refill_slots_4_way <= refill_push_payload_way;
        refill_slots_4_cmdSent <= 1'b0;
        refill_slots_4_priority <= 7'h7f;
        refill_slots_4_loaded <= 1'b0;
        refill_slots_4_loadedCounter <= 1'b0;
        refill_slots_4_victim <= refill_push_payload_victim;
        refill_slots_4_writebackHazards <= 8'h0;
      end else begin
        if(_zz_16) begin
          refill_slots_4_priority[0] <= 1'b0;
        end
        if(_zz_17) begin
          refill_slots_4_priority[1] <= 1'b0;
        end
        if(_zz_18) begin
          refill_slots_4_priority[2] <= 1'b0;
        end
        if(_zz_19) begin
          refill_slots_4_priority[3] <= 1'b0;
        end
        if(_zz_21) begin
          refill_slots_4_priority[4] <= 1'b0;
        end
        if(_zz_22) begin
          refill_slots_4_priority[5] <= 1'b0;
        end
        if(_zz_23) begin
          refill_slots_4_priority[6] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_dcache2_l750_5) begin
        refill_slots_5_address <= refill_push_payload_address;
        refill_slots_5_way <= refill_push_payload_way;
        refill_slots_5_cmdSent <= 1'b0;
        refill_slots_5_priority <= 7'h7f;
        refill_slots_5_loaded <= 1'b0;
        refill_slots_5_loadedCounter <= 1'b0;
        refill_slots_5_victim <= refill_push_payload_victim;
        refill_slots_5_writebackHazards <= 8'h0;
      end else begin
        if(_zz_16) begin
          refill_slots_5_priority[0] <= 1'b0;
        end
        if(_zz_17) begin
          refill_slots_5_priority[1] <= 1'b0;
        end
        if(_zz_18) begin
          refill_slots_5_priority[2] <= 1'b0;
        end
        if(_zz_19) begin
          refill_slots_5_priority[3] <= 1'b0;
        end
        if(_zz_20) begin
          refill_slots_5_priority[4] <= 1'b0;
        end
        if(_zz_22) begin
          refill_slots_5_priority[5] <= 1'b0;
        end
        if(_zz_23) begin
          refill_slots_5_priority[6] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_dcache2_l750_6) begin
        refill_slots_6_address <= refill_push_payload_address;
        refill_slots_6_way <= refill_push_payload_way;
        refill_slots_6_cmdSent <= 1'b0;
        refill_slots_6_priority <= 7'h7f;
        refill_slots_6_loaded <= 1'b0;
        refill_slots_6_loadedCounter <= 1'b0;
        refill_slots_6_victim <= refill_push_payload_victim;
        refill_slots_6_writebackHazards <= 8'h0;
      end else begin
        if(_zz_16) begin
          refill_slots_6_priority[0] <= 1'b0;
        end
        if(_zz_17) begin
          refill_slots_6_priority[1] <= 1'b0;
        end
        if(_zz_18) begin
          refill_slots_6_priority[2] <= 1'b0;
        end
        if(_zz_19) begin
          refill_slots_6_priority[3] <= 1'b0;
        end
        if(_zz_20) begin
          refill_slots_6_priority[4] <= 1'b0;
        end
        if(_zz_21) begin
          refill_slots_6_priority[5] <= 1'b0;
        end
        if(_zz_23) begin
          refill_slots_6_priority[6] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_dcache2_l750_7) begin
        refill_slots_7_address <= refill_push_payload_address;
        refill_slots_7_way <= refill_push_payload_way;
        refill_slots_7_cmdSent <= 1'b0;
        refill_slots_7_priority <= 7'h7f;
        refill_slots_7_loaded <= 1'b0;
        refill_slots_7_loadedCounter <= 1'b0;
        refill_slots_7_victim <= refill_push_payload_victim;
        refill_slots_7_writebackHazards <= 8'h0;
      end else begin
        if(_zz_16) begin
          refill_slots_7_priority[0] <= 1'b0;
        end
        if(_zz_17) begin
          refill_slots_7_priority[1] <= 1'b0;
        end
        if(_zz_18) begin
          refill_slots_7_priority[2] <= 1'b0;
        end
        if(_zz_19) begin
          refill_slots_7_priority[3] <= 1'b0;
        end
        if(_zz_20) begin
          refill_slots_7_priority[4] <= 1'b0;
        end
        if(_zz_21) begin
          refill_slots_7_priority[5] <= 1'b0;
        end
        if(_zz_22) begin
          refill_slots_7_priority[6] <= 1'b0;
        end
      end
    end
    if(refill_read_arbiter_oh[0]) begin
      refill_slots_0_writebackHazards <= refill_read_writebackHazards;
      if(when_dcache2_l791) begin
        refill_slots_0_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel) begin
      refill_slots_1_writebackHazards <= refill_read_writebackHazards;
      if(when_dcache2_l791_1) begin
        refill_slots_1_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel_1) begin
      refill_slots_2_writebackHazards <= refill_read_writebackHazards;
      if(when_dcache2_l791_2) begin
        refill_slots_2_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel_2) begin
      refill_slots_3_writebackHazards <= refill_read_writebackHazards;
      if(when_dcache2_l791_3) begin
        refill_slots_3_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel_3) begin
      refill_slots_4_writebackHazards <= refill_read_writebackHazards;
      if(when_dcache2_l791_4) begin
        refill_slots_4_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel_4) begin
      refill_slots_5_writebackHazards <= refill_read_writebackHazards;
      if(when_dcache2_l791_5) begin
        refill_slots_5_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel_5) begin
      refill_slots_6_writebackHazards <= refill_read_writebackHazards;
      if(when_dcache2_l791_6) begin
        refill_slots_6_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel_6) begin
      refill_slots_7_writebackHazards <= refill_read_writebackHazards;
      if(when_dcache2_l791_7) begin
        refill_slots_7_cmdSent <= 1'b1;
      end
    end
    if(io_mem_read_rsp_valid) begin
      if(when_dcache2_l834) begin
        case(io_mem_read_rsp_payload_id)
          3'b000 : begin
            refill_slots_0_loaded <= 1'b1;
          end
          3'b001 : begin
            refill_slots_1_loaded <= 1'b1;
          end
          3'b010 : begin
            refill_slots_2_loaded <= 1'b1;
          end
          3'b011 : begin
            refill_slots_3_loaded <= 1'b1;
          end
          3'b100 : begin
            refill_slots_4_loaded <= 1'b1;
          end
          3'b101 : begin
            refill_slots_5_loaded <= 1'b1;
          end
          3'b110 : begin
            refill_slots_6_loaded <= 1'b1;
          end
          default : begin
            refill_slots_7_loaded <= 1'b1;
          end
        endcase
      end
    end
    if(writeback_slots_0_fire) begin
      refill_slots_0_writebackHazards[0] <= 1'b0;
      refill_slots_1_writebackHazards[0] <= 1'b0;
      refill_slots_2_writebackHazards[0] <= 1'b0;
      refill_slots_3_writebackHazards[0] <= 1'b0;
      refill_slots_4_writebackHazards[0] <= 1'b0;
      refill_slots_5_writebackHazards[0] <= 1'b0;
      refill_slots_6_writebackHazards[0] <= 1'b0;
      refill_slots_7_writebackHazards[0] <= 1'b0;
    end
    if(writeback_slots_1_fire) begin
      refill_slots_0_writebackHazards[1] <= 1'b0;
      refill_slots_1_writebackHazards[1] <= 1'b0;
      refill_slots_2_writebackHazards[1] <= 1'b0;
      refill_slots_3_writebackHazards[1] <= 1'b0;
      refill_slots_4_writebackHazards[1] <= 1'b0;
      refill_slots_5_writebackHazards[1] <= 1'b0;
      refill_slots_6_writebackHazards[1] <= 1'b0;
      refill_slots_7_writebackHazards[1] <= 1'b0;
    end
    if(writeback_slots_2_fire) begin
      refill_slots_0_writebackHazards[2] <= 1'b0;
      refill_slots_1_writebackHazards[2] <= 1'b0;
      refill_slots_2_writebackHazards[2] <= 1'b0;
      refill_slots_3_writebackHazards[2] <= 1'b0;
      refill_slots_4_writebackHazards[2] <= 1'b0;
      refill_slots_5_writebackHazards[2] <= 1'b0;
      refill_slots_6_writebackHazards[2] <= 1'b0;
      refill_slots_7_writebackHazards[2] <= 1'b0;
    end
    if(writeback_slots_3_fire) begin
      refill_slots_0_writebackHazards[3] <= 1'b0;
      refill_slots_1_writebackHazards[3] <= 1'b0;
      refill_slots_2_writebackHazards[3] <= 1'b0;
      refill_slots_3_writebackHazards[3] <= 1'b0;
      refill_slots_4_writebackHazards[3] <= 1'b0;
      refill_slots_5_writebackHazards[3] <= 1'b0;
      refill_slots_6_writebackHazards[3] <= 1'b0;
      refill_slots_7_writebackHazards[3] <= 1'b0;
    end
    if(writeback_slots_4_fire) begin
      refill_slots_0_writebackHazards[4] <= 1'b0;
      refill_slots_1_writebackHazards[4] <= 1'b0;
      refill_slots_2_writebackHazards[4] <= 1'b0;
      refill_slots_3_writebackHazards[4] <= 1'b0;
      refill_slots_4_writebackHazards[4] <= 1'b0;
      refill_slots_5_writebackHazards[4] <= 1'b0;
      refill_slots_6_writebackHazards[4] <= 1'b0;
      refill_slots_7_writebackHazards[4] <= 1'b0;
    end
    if(writeback_slots_5_fire) begin
      refill_slots_0_writebackHazards[5] <= 1'b0;
      refill_slots_1_writebackHazards[5] <= 1'b0;
      refill_slots_2_writebackHazards[5] <= 1'b0;
      refill_slots_3_writebackHazards[5] <= 1'b0;
      refill_slots_4_writebackHazards[5] <= 1'b0;
      refill_slots_5_writebackHazards[5] <= 1'b0;
      refill_slots_6_writebackHazards[5] <= 1'b0;
      refill_slots_7_writebackHazards[5] <= 1'b0;
    end
    if(writeback_slots_6_fire) begin
      refill_slots_0_writebackHazards[6] <= 1'b0;
      refill_slots_1_writebackHazards[6] <= 1'b0;
      refill_slots_2_writebackHazards[6] <= 1'b0;
      refill_slots_3_writebackHazards[6] <= 1'b0;
      refill_slots_4_writebackHazards[6] <= 1'b0;
      refill_slots_5_writebackHazards[6] <= 1'b0;
      refill_slots_6_writebackHazards[6] <= 1'b0;
      refill_slots_7_writebackHazards[6] <= 1'b0;
    end
    if(writeback_slots_7_fire) begin
      refill_slots_0_writebackHazards[7] <= 1'b0;
      refill_slots_1_writebackHazards[7] <= 1'b0;
      refill_slots_2_writebackHazards[7] <= 1'b0;
      refill_slots_3_writebackHazards[7] <= 1'b0;
      refill_slots_4_writebackHazards[7] <= 1'b0;
      refill_slots_5_writebackHazards[7] <= 1'b0;
      refill_slots_6_writebackHazards[7] <= 1'b0;
      refill_slots_7_writebackHazards[7] <= 1'b0;
    end
    if(writeback_push_valid) begin
      if(when_dcache2_l897) begin
        writeback_slots_0_address <= writeback_push_payload_address;
        writeback_slots_0_way <= writeback_push_payload_way;
        writeback_slots_0_writeCmdDone <= 1'b0;
        writeback_slots_0_priority <= 7'h7f;
        writeback_slots_0_readCmdDone <= 1'b0;
        writeback_slots_0_readRspDone <= 1'b0;
        writeback_slots_0_victimBufferReady <= 1'b0;
      end else begin
        if(_zz_25) begin
          writeback_slots_0_priority[0] <= 1'b0;
        end
        if(_zz_26) begin
          writeback_slots_0_priority[1] <= 1'b0;
        end
        if(_zz_27) begin
          writeback_slots_0_priority[2] <= 1'b0;
        end
        if(_zz_28) begin
          writeback_slots_0_priority[3] <= 1'b0;
        end
        if(_zz_29) begin
          writeback_slots_0_priority[4] <= 1'b0;
        end
        if(_zz_30) begin
          writeback_slots_0_priority[5] <= 1'b0;
        end
        if(_zz_31) begin
          writeback_slots_0_priority[6] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_dcache2_l897_1) begin
        writeback_slots_1_address <= writeback_push_payload_address;
        writeback_slots_1_way <= writeback_push_payload_way;
        writeback_slots_1_writeCmdDone <= 1'b0;
        writeback_slots_1_priority <= 7'h7f;
        writeback_slots_1_readCmdDone <= 1'b0;
        writeback_slots_1_readRspDone <= 1'b0;
        writeback_slots_1_victimBufferReady <= 1'b0;
      end else begin
        if(_zz_24) begin
          writeback_slots_1_priority[0] <= 1'b0;
        end
        if(_zz_26) begin
          writeback_slots_1_priority[1] <= 1'b0;
        end
        if(_zz_27) begin
          writeback_slots_1_priority[2] <= 1'b0;
        end
        if(_zz_28) begin
          writeback_slots_1_priority[3] <= 1'b0;
        end
        if(_zz_29) begin
          writeback_slots_1_priority[4] <= 1'b0;
        end
        if(_zz_30) begin
          writeback_slots_1_priority[5] <= 1'b0;
        end
        if(_zz_31) begin
          writeback_slots_1_priority[6] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_dcache2_l897_2) begin
        writeback_slots_2_address <= writeback_push_payload_address;
        writeback_slots_2_way <= writeback_push_payload_way;
        writeback_slots_2_writeCmdDone <= 1'b0;
        writeback_slots_2_priority <= 7'h7f;
        writeback_slots_2_readCmdDone <= 1'b0;
        writeback_slots_2_readRspDone <= 1'b0;
        writeback_slots_2_victimBufferReady <= 1'b0;
      end else begin
        if(_zz_24) begin
          writeback_slots_2_priority[0] <= 1'b0;
        end
        if(_zz_25) begin
          writeback_slots_2_priority[1] <= 1'b0;
        end
        if(_zz_27) begin
          writeback_slots_2_priority[2] <= 1'b0;
        end
        if(_zz_28) begin
          writeback_slots_2_priority[3] <= 1'b0;
        end
        if(_zz_29) begin
          writeback_slots_2_priority[4] <= 1'b0;
        end
        if(_zz_30) begin
          writeback_slots_2_priority[5] <= 1'b0;
        end
        if(_zz_31) begin
          writeback_slots_2_priority[6] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_dcache2_l897_3) begin
        writeback_slots_3_address <= writeback_push_payload_address;
        writeback_slots_3_way <= writeback_push_payload_way;
        writeback_slots_3_writeCmdDone <= 1'b0;
        writeback_slots_3_priority <= 7'h7f;
        writeback_slots_3_readCmdDone <= 1'b0;
        writeback_slots_3_readRspDone <= 1'b0;
        writeback_slots_3_victimBufferReady <= 1'b0;
      end else begin
        if(_zz_24) begin
          writeback_slots_3_priority[0] <= 1'b0;
        end
        if(_zz_25) begin
          writeback_slots_3_priority[1] <= 1'b0;
        end
        if(_zz_26) begin
          writeback_slots_3_priority[2] <= 1'b0;
        end
        if(_zz_28) begin
          writeback_slots_3_priority[3] <= 1'b0;
        end
        if(_zz_29) begin
          writeback_slots_3_priority[4] <= 1'b0;
        end
        if(_zz_30) begin
          writeback_slots_3_priority[5] <= 1'b0;
        end
        if(_zz_31) begin
          writeback_slots_3_priority[6] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_dcache2_l897_4) begin
        writeback_slots_4_address <= writeback_push_payload_address;
        writeback_slots_4_way <= writeback_push_payload_way;
        writeback_slots_4_writeCmdDone <= 1'b0;
        writeback_slots_4_priority <= 7'h7f;
        writeback_slots_4_readCmdDone <= 1'b0;
        writeback_slots_4_readRspDone <= 1'b0;
        writeback_slots_4_victimBufferReady <= 1'b0;
      end else begin
        if(_zz_24) begin
          writeback_slots_4_priority[0] <= 1'b0;
        end
        if(_zz_25) begin
          writeback_slots_4_priority[1] <= 1'b0;
        end
        if(_zz_26) begin
          writeback_slots_4_priority[2] <= 1'b0;
        end
        if(_zz_27) begin
          writeback_slots_4_priority[3] <= 1'b0;
        end
        if(_zz_29) begin
          writeback_slots_4_priority[4] <= 1'b0;
        end
        if(_zz_30) begin
          writeback_slots_4_priority[5] <= 1'b0;
        end
        if(_zz_31) begin
          writeback_slots_4_priority[6] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_dcache2_l897_5) begin
        writeback_slots_5_address <= writeback_push_payload_address;
        writeback_slots_5_way <= writeback_push_payload_way;
        writeback_slots_5_writeCmdDone <= 1'b0;
        writeback_slots_5_priority <= 7'h7f;
        writeback_slots_5_readCmdDone <= 1'b0;
        writeback_slots_5_readRspDone <= 1'b0;
        writeback_slots_5_victimBufferReady <= 1'b0;
      end else begin
        if(_zz_24) begin
          writeback_slots_5_priority[0] <= 1'b0;
        end
        if(_zz_25) begin
          writeback_slots_5_priority[1] <= 1'b0;
        end
        if(_zz_26) begin
          writeback_slots_5_priority[2] <= 1'b0;
        end
        if(_zz_27) begin
          writeback_slots_5_priority[3] <= 1'b0;
        end
        if(_zz_28) begin
          writeback_slots_5_priority[4] <= 1'b0;
        end
        if(_zz_30) begin
          writeback_slots_5_priority[5] <= 1'b0;
        end
        if(_zz_31) begin
          writeback_slots_5_priority[6] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_dcache2_l897_6) begin
        writeback_slots_6_address <= writeback_push_payload_address;
        writeback_slots_6_way <= writeback_push_payload_way;
        writeback_slots_6_writeCmdDone <= 1'b0;
        writeback_slots_6_priority <= 7'h7f;
        writeback_slots_6_readCmdDone <= 1'b0;
        writeback_slots_6_readRspDone <= 1'b0;
        writeback_slots_6_victimBufferReady <= 1'b0;
      end else begin
        if(_zz_24) begin
          writeback_slots_6_priority[0] <= 1'b0;
        end
        if(_zz_25) begin
          writeback_slots_6_priority[1] <= 1'b0;
        end
        if(_zz_26) begin
          writeback_slots_6_priority[2] <= 1'b0;
        end
        if(_zz_27) begin
          writeback_slots_6_priority[3] <= 1'b0;
        end
        if(_zz_28) begin
          writeback_slots_6_priority[4] <= 1'b0;
        end
        if(_zz_29) begin
          writeback_slots_6_priority[5] <= 1'b0;
        end
        if(_zz_31) begin
          writeback_slots_6_priority[6] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_dcache2_l897_7) begin
        writeback_slots_7_address <= writeback_push_payload_address;
        writeback_slots_7_way <= writeback_push_payload_way;
        writeback_slots_7_writeCmdDone <= 1'b0;
        writeback_slots_7_priority <= 7'h7f;
        writeback_slots_7_readCmdDone <= 1'b0;
        writeback_slots_7_readRspDone <= 1'b0;
        writeback_slots_7_victimBufferReady <= 1'b0;
      end else begin
        if(_zz_24) begin
          writeback_slots_7_priority[0] <= 1'b0;
        end
        if(_zz_25) begin
          writeback_slots_7_priority[1] <= 1'b0;
        end
        if(_zz_26) begin
          writeback_slots_7_priority[2] <= 1'b0;
        end
        if(_zz_27) begin
          writeback_slots_7_priority[3] <= 1'b0;
        end
        if(_zz_28) begin
          writeback_slots_7_priority[4] <= 1'b0;
        end
        if(_zz_29) begin
          writeback_slots_7_priority[5] <= 1'b0;
        end
        if(_zz_30) begin
          writeback_slots_7_priority[6] <= 1'b0;
        end
      end
    end
    if(when_dcache2_l937) begin
      if(writeback_read_arbiter_oh[0]) begin
        writeback_slots_0_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel) begin
        writeback_slots_1_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel_1) begin
        writeback_slots_2_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel_2) begin
        writeback_slots_3_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel_3) begin
        writeback_slots_4_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel_4) begin
        writeback_slots_5_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel_5) begin
        writeback_slots_6_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel_6) begin
        writeback_slots_7_readCmdDone <= 1'b1;
      end
    end
    if(writeback_read_slotRead_valid) begin
      refill_slots_0_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_1_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_2_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_3_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_4_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_5_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_6_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_7_victim[writeback_read_slotRead_payload_id] <= 1'b0;
    end
    writeback_read_slotReadLast_payload_id <= writeback_read_slotRead_payload_id;
    writeback_read_slotReadLast_payload_last <= writeback_read_slotRead_payload_last;
    writeback_read_slotReadLast_payload_wordIndex <= writeback_read_slotRead_payload_wordIndex;
    writeback_read_slotReadLast_payload_way <= writeback_read_slotRead_payload_way;
    if(writeback_read_slotReadLast_valid) begin
      case(writeback_read_slotReadLast_payload_id)
        3'b000 : begin
          writeback_slots_0_victimBufferReady <= 1'b1;
        end
        3'b001 : begin
          writeback_slots_1_victimBufferReady <= 1'b1;
        end
        3'b010 : begin
          writeback_slots_2_victimBufferReady <= 1'b1;
        end
        3'b011 : begin
          writeback_slots_3_victimBufferReady <= 1'b1;
        end
        3'b100 : begin
          writeback_slots_4_victimBufferReady <= 1'b1;
        end
        3'b101 : begin
          writeback_slots_5_victimBufferReady <= 1'b1;
        end
        3'b110 : begin
          writeback_slots_6_victimBufferReady <= 1'b1;
        end
        default : begin
          writeback_slots_7_victimBufferReady <= 1'b1;
        end
      endcase
      if(writeback_read_slotReadLast_payload_last) begin
        case(writeback_read_slotReadLast_payload_id)
          3'b000 : begin
            writeback_slots_0_readRspDone <= 1'b1;
          end
          3'b001 : begin
            writeback_slots_1_readRspDone <= 1'b1;
          end
          3'b010 : begin
            writeback_slots_2_readRspDone <= 1'b1;
          end
          3'b011 : begin
            writeback_slots_3_readRspDone <= 1'b1;
          end
          3'b100 : begin
            writeback_slots_4_readRspDone <= 1'b1;
          end
          3'b101 : begin
            writeback_slots_5_readRspDone <= 1'b1;
          end
          3'b110 : begin
            writeback_slots_6_readRspDone <= 1'b1;
          end
          default : begin
            writeback_slots_7_readRspDone <= 1'b1;
          end
        endcase
      end
    end
    if(when_dcache2_l1020) begin
      if(writeback_write_arbiter_oh[0]) begin
        writeback_slots_0_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel) begin
        writeback_slots_1_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel_1) begin
        writeback_slots_2_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel_2) begin
        writeback_slots_3_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel_3) begin
        writeback_slots_4_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel_4) begin
        writeback_slots_5_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel_5) begin
        writeback_slots_6_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel_6) begin
        writeback_slots_7_writeCmdDone <= 1'b1;
      end
    end
    if(writeback_write_bufferRead_ready) begin
      writeback_write_bufferRead_rData_id <= writeback_write_bufferRead_payload_id;
      writeback_write_bufferRead_rData_address <= writeback_write_bufferRead_payload_address;
      writeback_write_bufferRead_rData_last <= writeback_write_bufferRead_payload_last;
    end
    load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION <= load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION;
    load_pipeline_stages_1_TRANSACTION_ID <= load_pipeline_stages_0_TRANSACTION_ID;
    load_pipeline_stages_1_WAYS_HAZARD <= load_pipeline_stages_0_WAYS_HAZARD;
    load_pipeline_stages_1_BANK_BUSY <= load_pipeline_stages_0_BANK_BUSY_overloaded;
    load_pipeline_stages_1_ADDRESS_POST_TRANSLATION <= load_pipeline_stages_0_ADDRESS_POST_TRANSLATION;
    load_pipeline_stages_1_ABORD <= load_pipeline_stages_0_ABORD;
    load_pipeline_stages_2_WAYS_HAZARD <= load_pipeline_stages_1_WAYS_HAZARD_overloaded;
    load_pipeline_stages_2_BANK_BUSY_REMAPPED <= load_pipeline_stages_1_BANK_BUSY_REMAPPED;
    load_pipeline_stages_2_BANKS_MUXES_0 <= load_pipeline_stages_1_BANKS_MUXES_0;
    load_pipeline_stages_2_BANKS_MUXES_1 <= load_pipeline_stages_1_BANKS_MUXES_1;
    load_pipeline_stages_2_WAYS_TAGS_0_loaded <= load_pipeline_stages_1_WAYS_TAGS_0_loaded;
    load_pipeline_stages_2_WAYS_TAGS_0_address <= load_pipeline_stages_1_WAYS_TAGS_0_address;
    load_pipeline_stages_2_WAYS_TAGS_0_fault <= load_pipeline_stages_1_WAYS_TAGS_0_fault;
    load_pipeline_stages_2_WAYS_TAGS_1_loaded <= load_pipeline_stages_1_WAYS_TAGS_1_loaded;
    load_pipeline_stages_2_WAYS_TAGS_1_address <= load_pipeline_stages_1_WAYS_TAGS_1_address;
    load_pipeline_stages_2_WAYS_TAGS_1_fault <= load_pipeline_stages_1_WAYS_TAGS_1_fault;
    load_pipeline_stages_2_WAYS_HITS <= load_pipeline_stages_1_WAYS_HITS;
    load_pipeline_stages_2_ADDRESS_POST_TRANSLATION <= load_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
    load_pipeline_stages_2_STATUS_0_dirty <= load_pipeline_stages_1_STATUS_overloaded_0_dirty;
    load_pipeline_stages_2_STATUS_1_dirty <= load_pipeline_stages_1_STATUS_overloaded_1_dirty;
    load_pipeline_stages_2_REFILL_HITS_EARLY <= load_pipeline_stages_1_REFILL_HITS_EARLY;
    load_pipeline_stages_2_ABORD <= load_pipeline_stages_1_ABORD;
    load_pipeline_stages_2_TRANSACTION_ID <= load_pipeline_stages_1_TRANSACTION_ID;
    store_pipeline_stages_1_ADDRESS_POST_TRANSLATION <= store_pipeline_stages_0_ADDRESS_POST_TRANSLATION;
    store_pipeline_stages_1_CPU_WORD <= store_pipeline_stages_0_CPU_WORD;
    store_pipeline_stages_1_CPU_MASK <= store_pipeline_stages_0_CPU_MASK;
    store_pipeline_stages_1_IO <= store_pipeline_stages_0_IO;
    store_pipeline_stages_1_FLUSH <= store_pipeline_stages_0_FLUSH;
    store_pipeline_stages_1_FLUSH_FREE <= store_pipeline_stages_0_FLUSH_FREE;
    store_pipeline_stages_1_PREFETCH <= store_pipeline_stages_0_PREFETCH;
    store_pipeline_stages_1_TRANSACTION_ID <= store_pipeline_stages_0_TRANSACTION_ID;
    store_pipeline_stages_1_WAYS_HAZARD <= store_pipeline_stages_0_WAYS_HAZARD;
    store_pipeline_stages_2_WAYS_HAZARD <= store_pipeline_stages_1_WAYS_HAZARD_overloaded;
    store_pipeline_stages_2_ADDRESS_POST_TRANSLATION <= store_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
    store_pipeline_stages_2_WAYS_TAGS_0_loaded <= store_pipeline_stages_1_WAYS_TAGS_0_loaded;
    store_pipeline_stages_2_WAYS_TAGS_0_address <= store_pipeline_stages_1_WAYS_TAGS_0_address;
    store_pipeline_stages_2_WAYS_TAGS_0_fault <= store_pipeline_stages_1_WAYS_TAGS_0_fault;
    store_pipeline_stages_2_WAYS_TAGS_1_loaded <= store_pipeline_stages_1_WAYS_TAGS_1_loaded;
    store_pipeline_stages_2_WAYS_TAGS_1_address <= store_pipeline_stages_1_WAYS_TAGS_1_address;
    store_pipeline_stages_2_WAYS_TAGS_1_fault <= store_pipeline_stages_1_WAYS_TAGS_1_fault;
    store_pipeline_stages_2_WAYS_HITS <= store_pipeline_stages_1_WAYS_HITS;
    store_pipeline_stages_2_WAYS_HIT <= store_pipeline_stages_1_WAYS_HIT;
    store_pipeline_stages_2_STATUS_0_dirty <= store_pipeline_stages_1_STATUS_overloaded_0_dirty;
    store_pipeline_stages_2_STATUS_1_dirty <= store_pipeline_stages_1_STATUS_overloaded_1_dirty;
    store_pipeline_stages_2_REFILL_HITS_EARLY <= store_pipeline_stages_1_REFILL_HITS_EARLY;
    store_pipeline_stages_2_FLUSH <= store_pipeline_stages_1_FLUSH;
    store_pipeline_stages_2_PREFETCH <= store_pipeline_stages_1_PREFETCH;
    store_pipeline_stages_2_IO <= store_pipeline_stages_1_IO;
    store_pipeline_stages_2_CPU_WORD <= store_pipeline_stages_1_CPU_WORD;
    store_pipeline_stages_2_CPU_MASK <= store_pipeline_stages_1_CPU_MASK;
    store_pipeline_stages_2_FLUSH_FREE <= store_pipeline_stages_1_FLUSH_FREE;
    store_pipeline_stages_2_TRANSACTION_ID <= store_pipeline_stages_1_TRANSACTION_ID;
  end

  always @(posedge clk) begin
    if(reset) begin
      status_writeLast_valid <= 1'b0;
      wayRandom_value <= 1'b0;
      invalidate_counter <= 5'h0;
      invalidate_done_regNext <= 1'b0;
      refill_slots_0_valid <= 1'b0;
      refill_slots_1_valid <= 1'b0;
      refill_slots_2_valid <= 1'b0;
      refill_slots_3_valid <= 1'b0;
      refill_slots_4_valid <= 1'b0;
      refill_slots_5_valid <= 1'b0;
      refill_slots_6_valid <= 1'b0;
      refill_slots_7_valid <= 1'b0;
      refill_read_arbiter_lock <= 8'h0;
      refill_read_wordIndex <= 3'b000;
      refill_read_hadError <= 1'b0;
      writeback_slots_0_valid <= 1'b0;
      writeback_slots_1_valid <= 1'b0;
      writeback_slots_2_valid <= 1'b0;
      writeback_slots_3_valid <= 1'b0;
      writeback_slots_4_valid <= 1'b0;
      writeback_slots_5_valid <= 1'b0;
      writeback_slots_6_valid <= 1'b0;
      writeback_slots_7_valid <= 1'b0;
      writeback_read_arbiter_lock <= 8'h0;
      writeback_read_wordIndex <= 3'b000;
      writeback_read_slotReadLast_valid <= 1'b0;
      writeback_write_arbiter_lock <= 8'h0;
      writeback_write_wordIndex <= 3'b000;
      writeback_write_bufferRead_rValid <= 1'b0;
      load_pipeline_stages_1_valid <= 1'b0;
      load_pipeline_stages_2_valid <= 1'b0;
      store_pipeline_stages_1_valid <= 1'b0;
      store_pipeline_stages_2_valid <= 1'b0;
    end else begin
      status_writeLast_valid <= status_write_valid;
      wayRandom_value <= wayRandom_valueNext;
      if(when_dcache2_l680) begin
        invalidate_counter <= (invalidate_counter + 5'h01);
      end
      invalidate_done_regNext <= invalidate_done;
      if(refill_slots_0_loadedDone) begin
        refill_slots_0_valid <= 1'b0;
      end
      if(refill_slots_1_loadedDone) begin
        refill_slots_1_valid <= 1'b0;
      end
      if(refill_slots_2_loadedDone) begin
        refill_slots_2_valid <= 1'b0;
      end
      if(refill_slots_3_loadedDone) begin
        refill_slots_3_valid <= 1'b0;
      end
      if(refill_slots_4_loadedDone) begin
        refill_slots_4_valid <= 1'b0;
      end
      if(refill_slots_5_loadedDone) begin
        refill_slots_5_valid <= 1'b0;
      end
      if(refill_slots_6_loadedDone) begin
        refill_slots_6_valid <= 1'b0;
      end
      if(refill_slots_7_loadedDone) begin
        refill_slots_7_valid <= 1'b0;
      end
      if(refill_push_valid) begin
        if(when_dcache2_l750) begin
          refill_slots_0_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_dcache2_l750_1) begin
          refill_slots_1_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_dcache2_l750_2) begin
          refill_slots_2_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_dcache2_l750_3) begin
          refill_slots_3_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_dcache2_l750_4) begin
          refill_slots_4_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_dcache2_l750_5) begin
          refill_slots_5_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_dcache2_l750_6) begin
          refill_slots_6_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_dcache2_l750_7) begin
          refill_slots_7_valid <= 1'b1;
        end
      end
      refill_read_arbiter_lock <= refill_read_arbiter_oh;
      if(when_dcache2_l779) begin
        refill_read_arbiter_lock <= 8'h0;
      end
      if(when_dcache2_l821) begin
        refill_read_hadError <= 1'b1;
      end
      if(io_mem_read_rsp_valid) begin
        if(refill_read_rspWithData) begin
          refill_read_wordIndex <= (refill_read_wordIndex + 3'b001);
        end
        if(when_dcache2_l834) begin
          refill_read_hadError <= 1'b0;
        end
      end
      if(writeback_slots_0_fire) begin
        writeback_slots_0_valid <= 1'b0;
      end
      if(writeback_slots_1_fire) begin
        writeback_slots_1_valid <= 1'b0;
      end
      if(writeback_slots_2_fire) begin
        writeback_slots_2_valid <= 1'b0;
      end
      if(writeback_slots_3_fire) begin
        writeback_slots_3_valid <= 1'b0;
      end
      if(writeback_slots_4_fire) begin
        writeback_slots_4_valid <= 1'b0;
      end
      if(writeback_slots_5_fire) begin
        writeback_slots_5_valid <= 1'b0;
      end
      if(writeback_slots_6_fire) begin
        writeback_slots_6_valid <= 1'b0;
      end
      if(writeback_slots_7_fire) begin
        writeback_slots_7_valid <= 1'b0;
      end
      if(writeback_push_valid) begin
        if(when_dcache2_l897) begin
          writeback_slots_0_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_dcache2_l897_1) begin
          writeback_slots_1_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_dcache2_l897_2) begin
          writeback_slots_2_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_dcache2_l897_3) begin
          writeback_slots_3_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_dcache2_l897_4) begin
          writeback_slots_4_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_dcache2_l897_5) begin
          writeback_slots_5_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_dcache2_l897_6) begin
          writeback_slots_6_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_dcache2_l897_7) begin
          writeback_slots_7_valid <= 1'b1;
        end
      end
      writeback_read_arbiter_lock <= writeback_read_arbiter_oh;
      writeback_read_wordIndex <= (writeback_read_wordIndex + _zz_writeback_read_wordIndex);
      if(when_dcache2_l937) begin
        writeback_read_arbiter_lock <= 8'h0;
      end
      writeback_read_slotReadLast_valid <= writeback_read_slotRead_valid;
      writeback_write_arbiter_lock <= writeback_write_arbiter_oh;
      writeback_write_wordIndex <= (writeback_write_wordIndex + _zz_writeback_write_wordIndex);
      if(when_dcache2_l1020) begin
        writeback_write_arbiter_lock <= 8'h0;
      end
      if(writeback_write_bufferRead_ready) begin
        writeback_write_bufferRead_rValid <= writeback_write_bufferRead_valid;
      end
      load_pipeline_stages_1_valid <= _zz_load_pipeline_stages_1_valid;
      load_pipeline_stages_2_valid <= _zz_load_pipeline_stages_2_valid;
      if(store_pipeline_stages_1_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // dcache2.scala:L1414
          `else
            if(!1'b0) begin
              $display("NOTE(dcache2.scala:1414):  [normal] [DCache] Store: Way 0 Tag read: loaded %x, address 0x%x, hit %x", store_pipeline_stages_1_WAYS_TAGS_0_loaded, store_pipeline_stages_1_WAYS_TAGS_0_address, _zz_35); // dcache2.scala:L1414
            end
          `endif
        `endif
      end
      if(store_pipeline_stages_1_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // dcache2.scala:L1414
          `else
            if(!1'b0) begin
              $display("NOTE(dcache2.scala:1414):  [normal] [DCache] Store: Way 1 Tag read: loaded %x, address 0x%x, hit %x", store_pipeline_stages_1_WAYS_TAGS_1_loaded, store_pipeline_stages_1_WAYS_TAGS_1_address, _zz_36); // dcache2.scala:L1414
            end
          `endif
        `endif
      end
      if(store_pipeline_stages_1_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // dcache2.scala:L1423
          `else
            if(!1'b0) begin
              $display("NOTE(dcache2.scala:1423):  [normal] [DCache] Store: Final hit decision: %x, ways hits: %x", _zz_37, _zz_38); // dcache2.scala:L1423
            end
          `endif
        `endif
      end
      if(store_ctrl_setDirty) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // dcache2.scala:L1604
          `else
            if(!1'b0) begin
              $display("NOTE(dcache2.scala:1604):  [normal] [DCache] STORE_SET_DIRTY: Address 0x%x, Line %x", _zz_39, _zz_40); // dcache2.scala:L1604
            end
          `endif
        `endif
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // dcache2.scala:L1605
          `else
            if(!1'b0) begin
              $display("NOTE(dcache2.scala:1605):  [normal] [DCache] STORE_SET_DIRTY: (controlStage )Address 0x%x, Line %x", store_pipeline_stages_2_ADDRESS_POST_TRANSLATION, _zz_41); // dcache2.scala:L1605
            end
          `endif
        `endif
      end
      if(store_pipeline_stages_2_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // dcache2.scala:L1626
          `else
            if(!1'b0) begin
              $display("NOTE(dcache2.scala:1626):  [normal] [DCache] Store: Control stage - WAYS_HIT: %x, MISS: %x, REDO: %x, IO: %x, FLUSH: %x, PREFETCH: %x", _zz_42, _zz_43, _zz_44, _zz_45, _zz_46, _zz_47); // dcache2.scala:L1626
            end
          `endif
        `endif
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // dcache2.scala:L1627
          `else
            if(!1'b0) begin
              $display("NOTE(dcache2.scala:1627):  [normal]   RefillHit: %x, LineBusy: %x, WaysHitHazard: %x, BankBusy: %x", store_ctrl_refillHit, store_ctrl_lineBusy, store_ctrl_waysHitHazard, store_ctrl_bankBusy); // dcache2.scala:L1627
            end
          `endif
        `endif
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // dcache2.scala:L1628
          `else
            if(!1'b0) begin
              $display("NOTE(dcache2.scala:1628):  [normal]   NeedFlush: %x, CanFlush: %x, StartFlush: %x", store_ctrl_needFlush, store_ctrl_canFlush, store_ctrl_startFlush); // dcache2.scala:L1628
            end
          `endif
        `endif
      end
      store_pipeline_stages_1_valid <= _zz_store_pipeline_stages_1_valid;
      store_pipeline_stages_2_valid <= _zz_store_pipeline_stages_2_valid;
    end
  end


endmodule

module SRAMController_1 (
  input  wire          io_axi_aw_valid,
  output reg           io_axi_aw_ready,
  input  wire [31:0]   io_axi_aw_payload_addr,
  input  wire [6:0]    io_axi_aw_payload_id,
  input  wire [7:0]    io_axi_aw_payload_len,
  input  wire [2:0]    io_axi_aw_payload_size,
  input  wire [1:0]    io_axi_aw_payload_burst,
  input  wire          io_axi_w_valid,
  output reg           io_axi_w_ready,
  input  wire [31:0]   io_axi_w_payload_data,
  input  wire [3:0]    io_axi_w_payload_strb,
  input  wire          io_axi_w_payload_last,
  output reg           io_axi_b_valid,
  input  wire          io_axi_b_ready,
  output reg  [6:0]    io_axi_b_payload_id,
  output reg  [1:0]    io_axi_b_payload_resp,
  input  wire          io_axi_ar_valid,
  output reg           io_axi_ar_ready,
  input  wire [31:0]   io_axi_ar_payload_addr,
  input  wire [6:0]    io_axi_ar_payload_id,
  input  wire [7:0]    io_axi_ar_payload_len,
  input  wire [2:0]    io_axi_ar_payload_size,
  input  wire [1:0]    io_axi_ar_payload_burst,
  output reg           io_axi_r_valid,
  input  wire          io_axi_r_ready,
  output reg  [31:0]   io_axi_r_payload_data,
  output reg  [6:0]    io_axi_r_payload_id,
  output reg  [1:0]    io_axi_r_payload_resp,
  output reg           io_axi_r_payload_last,
  input  wire [31:0]   io_ram_data_read,
  output wire [31:0]   io_ram_data_write,
  output wire          io_ram_data_writeEnable,
  output wire [19:0]   io_ram_addr,
  output wire [3:0]    io_ram_be_n,
  output wire          io_ram_ce_n,
  output wire          io_ram_oe_n,
  output wire          io_ram_we_n,
  input  wire          clk,
  input  wire          reset
);
  localparam fsm_BOOT = 4'd0;
  localparam fsm_IDLE = 4'd1;
  localparam fsm_VALIDATE = 4'd2;
  localparam fsm_WRITE_DATA_FETCH = 4'd3;
  localparam fsm_WRITE_EXECUTE = 4'd4;
  localparam fsm_WRITE_DEASSERT = 4'd5;
  localparam fsm_WRITE_FINALIZE = 4'd6;
  localparam fsm_WRITE_DATA_ERROR_CONSUME = 4'd7;
  localparam fsm_WRITE_RESPONSE = 4'd8;
  localparam fsm_READ_SETUP = 4'd9;
  localparam fsm_READ_WAIT = 4'd10;
  localparam fsm_READ_RESPONSE = 4'd11;
  localparam fsm_READ_RESPONSE_ERROR = 4'd12;

  wire       [7:0]    _zz_fsm_burst_count_remaining;
  wire       [17:0]   _zz_fsm_current_sram_addr;
  wire       [33:0]   _zz_fsm_current_sram_addr_1;
  wire       [33:0]   _zz_fsm_current_sram_addr_2;
  wire       [7:0]    _zz_fsm_burst_count_remaining_1;
  wire       [17:0]   _zz_fsm_current_sram_addr_3;
  wire       [33:0]   _zz_fsm_current_sram_addr_4;
  wire       [33:0]   _zz_fsm_current_sram_addr_5;
  wire       [19:0]   _zz_fsm_current_sram_addr_6;
  wire       [7:0]    _zz_fsm_current_sram_addr_7;
  wire       [7:0]    _zz_fsm_current_sram_addr_8;
  wire       [19:0]   _zz_fsm_next_sram_addr_prefetch;
  wire       [7:0]    _zz_fsm_next_sram_addr_prefetch_1;
  wire       [7:0]    _zz_fsm_next_sram_addr_prefetch_2;
  wire       [19:0]   _zz_fsm_current_sram_addr_9;
  wire       [7:0]    _zz_fsm_current_sram_addr_10;
  wire       [7:0]    _zz_fsm_current_sram_addr_11;
  wire       [3:0]    sram_be_n_inactive_value;
  (* mark_debug = "TRUE" *) reg        [19:0]   sram_addr_out_reg;
  (* mark_debug = "TRUE" *) reg        [31:0]   sram_data_out_reg;
  (* mark_debug = "TRUE" *) reg        [3:0]    sram_be_n_out_reg;
  (* mark_debug = "TRUE" *) reg                 sram_ce_n_out_reg;
  (* mark_debug = "TRUE" *) reg                 sram_oe_n_out_reg;
  (* mark_debug = "TRUE" *) reg                 sram_we_n_out_reg;
  (* mark_debug = "TRUE" *) reg                 sram_data_writeEnable_out_reg;
  (* mark_debug = "TRUE" *) reg        [31:0]   write_data_buffer;
  (* mark_debug = "TRUE" *) reg        [3:0]    write_strb_buffer;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  (* mark_debug = "TRUE" *) reg        [31:0]   fsm_ar_cmd_reg_addr;
  (* mark_debug = "TRUE" *) reg        [6:0]    fsm_ar_cmd_reg_id;
  (* mark_debug = "TRUE" *) reg        [7:0]    fsm_ar_cmd_reg_len;
  (* mark_debug = "TRUE" *) reg        [2:0]    fsm_ar_cmd_reg_size;
  (* mark_debug = "TRUE" *) reg        [1:0]    fsm_ar_cmd_reg_burst;
  (* mark_debug = "TRUE" *) reg        [31:0]   fsm_aw_cmd_reg_addr;
  (* mark_debug = "TRUE" *) reg        [6:0]    fsm_aw_cmd_reg_id;
  (* mark_debug = "TRUE" *) reg        [7:0]    fsm_aw_cmd_reg_len;
  (* mark_debug = "TRUE" *) reg        [2:0]    fsm_aw_cmd_reg_size;
  (* mark_debug = "TRUE" *) reg        [1:0]    fsm_aw_cmd_reg_burst;
  (* mark_debug = "TRUE" *) reg        [8:0]    fsm_burst_count_remaining;
  (* mark_debug = "TRUE" *) reg        [19:0]   fsm_current_sram_addr;
  (* mark_debug = "TRUE" *) reg        [31:0]   fsm_read_data_buffer;
  reg        [1:0]    fsm_read_wait_counter;
  reg        [1:0]    fsm_write_wait_counter;
  (* MARK_DEBUG = "TRUE" *) reg                 fsm_transaction_error_occurred;
  reg                 fsm_read_priority;
  reg        [19:0]   fsm_next_sram_addr_prefetch;
  reg                 fsm_addr_prefetch_valid;
  (* MARK_DEBUG = "TRUE" *) reg        [3:0]    fsm_stateReg;
  reg        [3:0]    fsm_stateNext;
  wire                when_SRAMController_l293;
  (* mark_debug = "true" *) wire                io_axi_aw_fire;
  (* mark_debug = "true" *) wire                io_axi_ar_fire;
  (* mark_debug = "true" *) wire                io_axi_w_fire;
  wire                when_SRAMController_l454;
  wire                when_SRAMController_l473;
  wire                when_SRAMController_l490;
  wire                when_SRAMController_l523;
  wire                when_SRAMController_l625;
  wire                when_SRAMController_l634;
  wire                when_SRAMController_l664;
  (* mark_debug = "true" *) wire                io_axi_r_fire;
  wire                when_SRAMController_l713;
  wire                fsm_onExit_BOOT;
  wire                fsm_onExit_IDLE;
  wire                fsm_onExit_VALIDATE;
  wire                fsm_onExit_WRITE_DATA_FETCH;
  wire                fsm_onExit_WRITE_EXECUTE;
  wire                fsm_onExit_WRITE_DEASSERT;
  wire                fsm_onExit_WRITE_FINALIZE;
  wire                fsm_onExit_WRITE_DATA_ERROR_CONSUME;
  wire                fsm_onExit_WRITE_RESPONSE;
  wire                fsm_onExit_READ_SETUP;
  wire                fsm_onExit_READ_WAIT;
  wire                fsm_onExit_READ_RESPONSE;
  wire                fsm_onExit_READ_RESPONSE_ERROR;
  wire                fsm_onEntry_BOOT;
  wire                fsm_onEntry_IDLE;
  wire                fsm_onEntry_VALIDATE;
  wire                fsm_onEntry_WRITE_DATA_FETCH;
  wire                fsm_onEntry_WRITE_EXECUTE;
  wire                fsm_onEntry_WRITE_DEASSERT;
  wire                fsm_onEntry_WRITE_FINALIZE;
  wire                fsm_onEntry_WRITE_DATA_ERROR_CONSUME;
  wire                fsm_onEntry_WRITE_RESPONSE;
  wire                fsm_onEntry_READ_SETUP;
  wire                fsm_onEntry_READ_WAIT;
  wire                fsm_onEntry_READ_RESPONSE;
  wire                fsm_onEntry_READ_RESPONSE_ERROR;
  (* mark_debug = "true" *) wire                io_axi_b_fire;
  reg                 sram_ce_n_out_reg_prev;
  reg                 sram_we_n_out_reg_prev;
  wire                when_SRAMController_l749;
  wire                when_SRAMController_l750;
  `ifndef SYNTHESIS
  reg [191:0] fsm_stateReg_string;
  reg [191:0] fsm_stateNext_string;
  `endif


  assign _zz_fsm_burst_count_remaining = (io_axi_aw_payload_len + 8'h01);
  assign _zz_fsm_current_sram_addr = (_zz_fsm_current_sram_addr_1[19 : 0] >>> 2'd2);
  assign _zz_fsm_current_sram_addr_1 = (_zz_fsm_current_sram_addr_2 - 34'h080400000);
  assign _zz_fsm_current_sram_addr_2 = {2'd0, io_axi_aw_payload_addr};
  assign _zz_fsm_burst_count_remaining_1 = (io_axi_ar_payload_len + 8'h01);
  assign _zz_fsm_current_sram_addr_3 = (_zz_fsm_current_sram_addr_4[19 : 0] >>> 2'd2);
  assign _zz_fsm_current_sram_addr_4 = (_zz_fsm_current_sram_addr_5 - 34'h080400000);
  assign _zz_fsm_current_sram_addr_5 = {2'd0, io_axi_ar_payload_addr};
  assign _zz_fsm_current_sram_addr_7 = (_zz_fsm_current_sram_addr_8 / 3'b100);
  assign _zz_fsm_current_sram_addr_6 = {12'd0, _zz_fsm_current_sram_addr_7};
  assign _zz_fsm_current_sram_addr_8 = ({7'd0,1'b1} <<< fsm_aw_cmd_reg_size);
  assign _zz_fsm_next_sram_addr_prefetch_1 = (_zz_fsm_next_sram_addr_prefetch_2 / 3'b100);
  assign _zz_fsm_next_sram_addr_prefetch = {12'd0, _zz_fsm_next_sram_addr_prefetch_1};
  assign _zz_fsm_next_sram_addr_prefetch_2 = ({7'd0,1'b1} <<< fsm_ar_cmd_reg_size);
  assign _zz_fsm_current_sram_addr_10 = (_zz_fsm_current_sram_addr_11 / 3'b100);
  assign _zz_fsm_current_sram_addr_9 = {12'd0, _zz_fsm_current_sram_addr_10};
  assign _zz_fsm_current_sram_addr_11 = ({7'd0,1'b1} <<< fsm_ar_cmd_reg_size);
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_BOOT : fsm_stateReg_string = "BOOT                    ";
      fsm_IDLE : fsm_stateReg_string = "IDLE                    ";
      fsm_VALIDATE : fsm_stateReg_string = "VALIDATE                ";
      fsm_WRITE_DATA_FETCH : fsm_stateReg_string = "WRITE_DATA_FETCH        ";
      fsm_WRITE_EXECUTE : fsm_stateReg_string = "WRITE_EXECUTE           ";
      fsm_WRITE_DEASSERT : fsm_stateReg_string = "WRITE_DEASSERT          ";
      fsm_WRITE_FINALIZE : fsm_stateReg_string = "WRITE_FINALIZE          ";
      fsm_WRITE_DATA_ERROR_CONSUME : fsm_stateReg_string = "WRITE_DATA_ERROR_CONSUME";
      fsm_WRITE_RESPONSE : fsm_stateReg_string = "WRITE_RESPONSE          ";
      fsm_READ_SETUP : fsm_stateReg_string = "READ_SETUP              ";
      fsm_READ_WAIT : fsm_stateReg_string = "READ_WAIT               ";
      fsm_READ_RESPONSE : fsm_stateReg_string = "READ_RESPONSE           ";
      fsm_READ_RESPONSE_ERROR : fsm_stateReg_string = "READ_RESPONSE_ERROR     ";
      default : fsm_stateReg_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_BOOT : fsm_stateNext_string = "BOOT                    ";
      fsm_IDLE : fsm_stateNext_string = "IDLE                    ";
      fsm_VALIDATE : fsm_stateNext_string = "VALIDATE                ";
      fsm_WRITE_DATA_FETCH : fsm_stateNext_string = "WRITE_DATA_FETCH        ";
      fsm_WRITE_EXECUTE : fsm_stateNext_string = "WRITE_EXECUTE           ";
      fsm_WRITE_DEASSERT : fsm_stateNext_string = "WRITE_DEASSERT          ";
      fsm_WRITE_FINALIZE : fsm_stateNext_string = "WRITE_FINALIZE          ";
      fsm_WRITE_DATA_ERROR_CONSUME : fsm_stateNext_string = "WRITE_DATA_ERROR_CONSUME";
      fsm_WRITE_RESPONSE : fsm_stateNext_string = "WRITE_RESPONSE          ";
      fsm_READ_SETUP : fsm_stateNext_string = "READ_SETUP              ";
      fsm_READ_WAIT : fsm_stateNext_string = "READ_WAIT               ";
      fsm_READ_RESPONSE : fsm_stateNext_string = "READ_RESPONSE           ";
      fsm_READ_RESPONSE_ERROR : fsm_stateNext_string = "READ_RESPONSE_ERROR     ";
      default : fsm_stateNext_string = "????????????????????????";
    endcase
  end
  `endif

  always @(*) begin
    io_axi_aw_ready = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
        io_axi_aw_ready = 1'b0;
        if(when_SRAMController_l293) begin
          io_axi_aw_ready = (! fsm_read_priority);
        end else begin
          io_axi_aw_ready = io_axi_aw_valid;
        end
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        io_axi_aw_ready = 1'b0;
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_ar_ready = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
        io_axi_ar_ready = 1'b0;
        if(when_SRAMController_l293) begin
          io_axi_ar_ready = fsm_read_priority;
        end else begin
          io_axi_ar_ready = io_axi_ar_valid;
        end
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        io_axi_ar_ready = 1'b0;
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_w_ready = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
        io_axi_w_ready = 1'b0;
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
        io_axi_w_ready = 1'b1;
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        io_axi_w_ready = 1'b1;
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_b_valid = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
        io_axi_b_valid = 1'b1;
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_valid = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_valid = 1'b1;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_b_payload_id = 7'h0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
        io_axi_b_payload_id = fsm_aw_cmd_reg_id;
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_b_payload_resp = 2'b00;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
        io_axi_b_payload_resp = (fsm_transaction_error_occurred ? 2'b10 : 2'b00);
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_payload_id = 7'h0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_payload_id = fsm_ar_cmd_reg_id;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_payload_id = fsm_ar_cmd_reg_id;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_payload_data = 32'h0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_payload_data = fsm_read_data_buffer;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_payload_data = 32'h0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_payload_resp = 2'b00;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_payload_resp = 2'b00;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_payload_resp = 2'b10;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_payload_last = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_payload_last = when_SRAMController_l664;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_payload_last = when_SRAMController_l713;
      end
      default : begin
      end
    endcase
  end

  assign sram_be_n_inactive_value = 4'b1111;
  assign io_ram_addr = sram_addr_out_reg;
  assign io_ram_ce_n = sram_ce_n_out_reg;
  assign io_ram_oe_n = sram_oe_n_out_reg;
  assign io_ram_we_n = sram_we_n_out_reg;
  assign io_ram_be_n = sram_be_n_out_reg;
  assign io_ram_data_write = sram_data_out_reg;
  assign io_ram_data_writeEnable = sram_data_writeEnable_out_reg;
  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_IDLE : begin
        if(io_axi_aw_fire) begin
          fsm_stateNext = fsm_WRITE_DATA_FETCH;
        end
        if(io_axi_ar_fire) begin
          fsm_stateNext = fsm_READ_SETUP;
        end
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
        if(io_axi_w_fire) begin
          fsm_stateNext = fsm_WRITE_EXECUTE;
        end
      end
      fsm_WRITE_EXECUTE : begin
        if(when_SRAMController_l454) begin
          fsm_stateNext = fsm_WRITE_DEASSERT;
        end
      end
      fsm_WRITE_DEASSERT : begin
        if(when_SRAMController_l473) begin
          fsm_stateNext = fsm_WRITE_FINALIZE;
        end
      end
      fsm_WRITE_FINALIZE : begin
        if(when_SRAMController_l490) begin
          fsm_stateNext = fsm_WRITE_RESPONSE;
        end else begin
          fsm_stateNext = fsm_WRITE_DATA_FETCH;
        end
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        if(io_axi_w_fire) begin
          if(when_SRAMController_l523) begin
            fsm_stateNext = fsm_WRITE_RESPONSE;
          end
        end
      end
      fsm_WRITE_RESPONSE : begin
        if(io_axi_b_ready) begin
          fsm_stateNext = fsm_IDLE;
        end
      end
      fsm_READ_SETUP : begin
        fsm_stateNext = fsm_READ_WAIT;
      end
      fsm_READ_WAIT : begin
        if(when_SRAMController_l634) begin
          fsm_stateNext = fsm_READ_RESPONSE;
        end
      end
      fsm_READ_RESPONSE : begin
        if(io_axi_r_fire) begin
          if(when_SRAMController_l664) begin
            fsm_stateNext = fsm_IDLE;
          end else begin
            fsm_stateNext = fsm_READ_SETUP;
          end
        end
      end
      fsm_READ_RESPONSE_ERROR : begin
        if(io_axi_r_fire) begin
          if(when_SRAMController_l713) begin
            fsm_stateNext = fsm_IDLE;
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_IDLE;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_BOOT;
    end
  end

  assign when_SRAMController_l293 = (io_axi_aw_valid && io_axi_ar_valid);
  assign io_axi_aw_fire = (io_axi_aw_valid && io_axi_aw_ready);
  assign io_axi_ar_fire = (io_axi_ar_valid && io_axi_ar_ready);
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign when_SRAMController_l454 = (fsm_write_wait_counter == 2'b11);
  assign when_SRAMController_l473 = 1'b1;
  assign when_SRAMController_l490 = (fsm_burst_count_remaining == 9'h0);
  assign when_SRAMController_l523 = (fsm_burst_count_remaining == 9'h001);
  assign when_SRAMController_l625 = (((fsm_read_wait_counter == 2'b10) && (9'h001 < fsm_burst_count_remaining)) && (! fsm_addr_prefetch_valid));
  assign when_SRAMController_l634 = (fsm_read_wait_counter == 2'b11);
  assign when_SRAMController_l664 = (fsm_burst_count_remaining == 9'h001);
  assign io_axi_r_fire = (io_axi_r_valid && io_axi_r_ready);
  assign when_SRAMController_l713 = (fsm_burst_count_remaining == 9'h001);
  assign fsm_onExit_BOOT = ((fsm_stateNext != fsm_BOOT) && (fsm_stateReg == fsm_BOOT));
  assign fsm_onExit_IDLE = ((fsm_stateNext != fsm_IDLE) && (fsm_stateReg == fsm_IDLE));
  assign fsm_onExit_VALIDATE = ((fsm_stateNext != fsm_VALIDATE) && (fsm_stateReg == fsm_VALIDATE));
  assign fsm_onExit_WRITE_DATA_FETCH = ((fsm_stateNext != fsm_WRITE_DATA_FETCH) && (fsm_stateReg == fsm_WRITE_DATA_FETCH));
  assign fsm_onExit_WRITE_EXECUTE = ((fsm_stateNext != fsm_WRITE_EXECUTE) && (fsm_stateReg == fsm_WRITE_EXECUTE));
  assign fsm_onExit_WRITE_DEASSERT = ((fsm_stateNext != fsm_WRITE_DEASSERT) && (fsm_stateReg == fsm_WRITE_DEASSERT));
  assign fsm_onExit_WRITE_FINALIZE = ((fsm_stateNext != fsm_WRITE_FINALIZE) && (fsm_stateReg == fsm_WRITE_FINALIZE));
  assign fsm_onExit_WRITE_DATA_ERROR_CONSUME = ((fsm_stateNext != fsm_WRITE_DATA_ERROR_CONSUME) && (fsm_stateReg == fsm_WRITE_DATA_ERROR_CONSUME));
  assign fsm_onExit_WRITE_RESPONSE = ((fsm_stateNext != fsm_WRITE_RESPONSE) && (fsm_stateReg == fsm_WRITE_RESPONSE));
  assign fsm_onExit_READ_SETUP = ((fsm_stateNext != fsm_READ_SETUP) && (fsm_stateReg == fsm_READ_SETUP));
  assign fsm_onExit_READ_WAIT = ((fsm_stateNext != fsm_READ_WAIT) && (fsm_stateReg == fsm_READ_WAIT));
  assign fsm_onExit_READ_RESPONSE = ((fsm_stateNext != fsm_READ_RESPONSE) && (fsm_stateReg == fsm_READ_RESPONSE));
  assign fsm_onExit_READ_RESPONSE_ERROR = ((fsm_stateNext != fsm_READ_RESPONSE_ERROR) && (fsm_stateReg == fsm_READ_RESPONSE_ERROR));
  assign fsm_onEntry_BOOT = ((fsm_stateNext == fsm_BOOT) && (fsm_stateReg != fsm_BOOT));
  assign fsm_onEntry_IDLE = ((fsm_stateNext == fsm_IDLE) && (fsm_stateReg != fsm_IDLE));
  assign fsm_onEntry_VALIDATE = ((fsm_stateNext == fsm_VALIDATE) && (fsm_stateReg != fsm_VALIDATE));
  assign fsm_onEntry_WRITE_DATA_FETCH = ((fsm_stateNext == fsm_WRITE_DATA_FETCH) && (fsm_stateReg != fsm_WRITE_DATA_FETCH));
  assign fsm_onEntry_WRITE_EXECUTE = ((fsm_stateNext == fsm_WRITE_EXECUTE) && (fsm_stateReg != fsm_WRITE_EXECUTE));
  assign fsm_onEntry_WRITE_DEASSERT = ((fsm_stateNext == fsm_WRITE_DEASSERT) && (fsm_stateReg != fsm_WRITE_DEASSERT));
  assign fsm_onEntry_WRITE_FINALIZE = ((fsm_stateNext == fsm_WRITE_FINALIZE) && (fsm_stateReg != fsm_WRITE_FINALIZE));
  assign fsm_onEntry_WRITE_DATA_ERROR_CONSUME = ((fsm_stateNext == fsm_WRITE_DATA_ERROR_CONSUME) && (fsm_stateReg != fsm_WRITE_DATA_ERROR_CONSUME));
  assign fsm_onEntry_WRITE_RESPONSE = ((fsm_stateNext == fsm_WRITE_RESPONSE) && (fsm_stateReg != fsm_WRITE_RESPONSE));
  assign fsm_onEntry_READ_SETUP = ((fsm_stateNext == fsm_READ_SETUP) && (fsm_stateReg != fsm_READ_SETUP));
  assign fsm_onEntry_READ_WAIT = ((fsm_stateNext == fsm_READ_WAIT) && (fsm_stateReg != fsm_READ_WAIT));
  assign fsm_onEntry_READ_RESPONSE = ((fsm_stateNext == fsm_READ_RESPONSE) && (fsm_stateReg != fsm_READ_RESPONSE));
  assign fsm_onEntry_READ_RESPONSE_ERROR = ((fsm_stateNext == fsm_READ_RESPONSE_ERROR) && (fsm_stateReg != fsm_READ_RESPONSE_ERROR));
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  assign when_SRAMController_l749 = ((sram_ce_n_out_reg_prev == 1'b0) && (sram_we_n_out_reg_prev == 1'b0));
  assign when_SRAMController_l750 = ((sram_ce_n_out_reg == 1'b1) && (sram_we_n_out_reg == 1'b1));
  always @(posedge clk) begin
    if(reset) begin
      sram_addr_out_reg <= 20'h0;
      sram_data_out_reg <= 32'h0;
      sram_be_n_out_reg <= sram_be_n_inactive_value;
      sram_ce_n_out_reg <= 1'b1;
      sram_oe_n_out_reg <= 1'b1;
      sram_we_n_out_reg <= 1'b1;
      sram_data_writeEnable_out_reg <= 1'b0;
      fsm_transaction_error_occurred <= 1'b0;
      fsm_read_priority <= 1'b0;
      fsm_addr_prefetch_valid <= 1'b0;
      fsm_stateReg <= fsm_BOOT;
      sram_ce_n_out_reg_prev <= 1'b1;
      sram_we_n_out_reg_prev <= 1'b1;
    end else begin
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_IDLE : begin
          fsm_transaction_error_occurred <= 1'b0;
          fsm_addr_prefetch_valid <= 1'b0;
          if(io_axi_aw_fire) begin
            fsm_read_priority <= (! fsm_read_priority);
            fsm_transaction_error_occurred <= 1'b0;
          end
          if(io_axi_ar_fire) begin
            fsm_read_priority <= (! fsm_read_priority);
            fsm_transaction_error_occurred <= 1'b0;
          end
        end
        fsm_VALIDATE : begin
        end
        fsm_WRITE_DATA_FETCH : begin
        end
        fsm_WRITE_EXECUTE : begin
        end
        fsm_WRITE_DEASSERT : begin
        end
        fsm_WRITE_FINALIZE : begin
        end
        fsm_WRITE_DATA_ERROR_CONSUME : begin
        end
        fsm_WRITE_RESPONSE : begin
        end
        fsm_READ_SETUP : begin
          fsm_addr_prefetch_valid <= 1'b0;
          sram_ce_n_out_reg <= 1'b0;
          sram_oe_n_out_reg <= 1'b0;
          sram_we_n_out_reg <= 1'b1;
          sram_data_writeEnable_out_reg <= 1'b0;
          sram_addr_out_reg <= fsm_current_sram_addr;
          sram_be_n_out_reg <= 4'b0000;
        end
        fsm_READ_WAIT : begin
          if(when_SRAMController_l625) begin
            fsm_addr_prefetch_valid <= 1'b1;
          end
        end
        fsm_READ_RESPONSE : begin
          if(io_axi_r_fire) begin
            if(!when_SRAMController_l664) begin
              if(fsm_addr_prefetch_valid) begin
                fsm_addr_prefetch_valid <= 1'b0;
              end
            end
          end
        end
        fsm_READ_RESPONSE_ERROR : begin
        end
        default : begin
        end
      endcase
      if(fsm_onExit_READ_RESPONSE) begin
        sram_oe_n_out_reg <= 1'b1;
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= sram_be_n_inactive_value;
        sram_addr_out_reg <= 20'h0;
      end
      if(fsm_onEntry_IDLE) begin
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
        sram_oe_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= sram_be_n_inactive_value;
        sram_addr_out_reg <= 20'h0;
      end
      if(fsm_onEntry_WRITE_DATA_FETCH) begin
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
      end
      if(fsm_onEntry_WRITE_EXECUTE) begin
        sram_addr_out_reg <= fsm_current_sram_addr;
        sram_data_out_reg <= io_axi_w_payload_data;
        sram_data_writeEnable_out_reg <= 1'b1;
        sram_be_n_out_reg <= (~ io_axi_w_payload_strb);
        sram_ce_n_out_reg <= 1'b0;
        sram_oe_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b0;
      end
      if(fsm_onEntry_WRITE_DEASSERT) begin
        sram_we_n_out_reg <= 1'b1;
      end
      if(fsm_onEntry_WRITE_FINALIZE) begin
        sram_ce_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
      end
      if(fsm_onEntry_WRITE_DATA_ERROR_CONSUME) begin
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
        sram_oe_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= sram_be_n_inactive_value;
        sram_addr_out_reg <= 20'h0;
      end
      if(fsm_onEntry_WRITE_RESPONSE) begin
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
        sram_oe_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= sram_be_n_inactive_value;
        sram_addr_out_reg <= 20'h0;
      end
      if(fsm_onEntry_READ_SETUP) begin
        sram_ce_n_out_reg <= 1'b0;
        sram_oe_n_out_reg <= 1'b0;
        sram_we_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_addr_out_reg <= fsm_current_sram_addr;
        sram_be_n_out_reg <= 4'b0000;
      end
      if(fsm_onEntry_READ_WAIT) begin
        sram_ce_n_out_reg <= 1'b0;
        sram_oe_n_out_reg <= 1'b0;
        sram_we_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= 4'b0000;
      end
      sram_ce_n_out_reg_prev <= sram_ce_n_out_reg;
      sram_we_n_out_reg_prev <= sram_we_n_out_reg;
      if(when_SRAMController_l749) begin
        if(when_SRAMController_l750) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // SRAMController.scala:L751
            `else
              if(!1'b0) begin
                $display("FAILURE This is a bug."); // SRAMController.scala:L751
                $finish;
              end
            `endif
          `endif
        end
      end
    end
  end

  always @(posedge clk) begin
    case(fsm_stateReg)
      fsm_IDLE : begin
        if(io_axi_aw_fire) begin
          fsm_aw_cmd_reg_addr <= io_axi_aw_payload_addr;
          fsm_aw_cmd_reg_id <= io_axi_aw_payload_id;
          fsm_aw_cmd_reg_len <= io_axi_aw_payload_len;
          fsm_aw_cmd_reg_size <= io_axi_aw_payload_size;
          fsm_aw_cmd_reg_burst <= io_axi_aw_payload_burst;
          fsm_burst_count_remaining <= {1'd0, _zz_fsm_burst_count_remaining};
          fsm_current_sram_addr <= {2'd0, _zz_fsm_current_sram_addr};
        end
        if(io_axi_ar_fire) begin
          fsm_ar_cmd_reg_addr <= io_axi_ar_payload_addr;
          fsm_ar_cmd_reg_id <= io_axi_ar_payload_id;
          fsm_ar_cmd_reg_len <= io_axi_ar_payload_len;
          fsm_ar_cmd_reg_size <= io_axi_ar_payload_size;
          fsm_ar_cmd_reg_burst <= io_axi_ar_payload_burst;
          fsm_burst_count_remaining <= {1'd0, _zz_fsm_burst_count_remaining_1};
          fsm_current_sram_addr <= {2'd0, _zz_fsm_current_sram_addr_3};
          fsm_read_wait_counter <= 2'b00;
        end
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
        if(when_SRAMController_l454) begin
          fsm_burst_count_remaining <= (fsm_burst_count_remaining - 9'h001);
        end else begin
          fsm_write_wait_counter <= (fsm_write_wait_counter + 2'b01);
        end
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
        if(!when_SRAMController_l490) begin
          fsm_current_sram_addr <= (fsm_current_sram_addr + _zz_fsm_current_sram_addr_6);
        end
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        if(io_axi_w_fire) begin
          fsm_burst_count_remaining <= (fsm_burst_count_remaining - 9'h001);
        end
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
        fsm_read_wait_counter <= 2'b00;
      end
      fsm_READ_WAIT : begin
        if(when_SRAMController_l625) begin
          fsm_next_sram_addr_prefetch <= (fsm_current_sram_addr + _zz_fsm_next_sram_addr_prefetch);
        end
        if(when_SRAMController_l634) begin
          fsm_read_data_buffer <= io_ram_data_read;
        end else begin
          fsm_read_wait_counter <= (fsm_read_wait_counter + 2'b01);
        end
      end
      fsm_READ_RESPONSE : begin
        if(io_axi_r_fire) begin
          fsm_burst_count_remaining <= (fsm_burst_count_remaining - 9'h001);
          if(!when_SRAMController_l664) begin
            if(fsm_addr_prefetch_valid) begin
              fsm_current_sram_addr <= fsm_next_sram_addr_prefetch;
            end else begin
              fsm_current_sram_addr <= (fsm_current_sram_addr + _zz_fsm_current_sram_addr_9);
            end
          end
        end
      end
      fsm_READ_RESPONSE_ERROR : begin
        if(io_axi_r_fire) begin
          fsm_burst_count_remaining <= (fsm_burst_count_remaining - 9'h001);
        end
      end
      default : begin
      end
    endcase
    if(fsm_onEntry_WRITE_EXECUTE) begin
      fsm_write_wait_counter <= 2'b00;
    end
  end


endmodule

module SRAMController (
  input  wire          io_axi_aw_valid,
  output reg           io_axi_aw_ready,
  input  wire [31:0]   io_axi_aw_payload_addr,
  input  wire [6:0]    io_axi_aw_payload_id,
  input  wire [7:0]    io_axi_aw_payload_len,
  input  wire [2:0]    io_axi_aw_payload_size,
  input  wire [1:0]    io_axi_aw_payload_burst,
  input  wire          io_axi_w_valid,
  output reg           io_axi_w_ready,
  input  wire [31:0]   io_axi_w_payload_data,
  input  wire [3:0]    io_axi_w_payload_strb,
  input  wire          io_axi_w_payload_last,
  output reg           io_axi_b_valid,
  input  wire          io_axi_b_ready,
  output reg  [6:0]    io_axi_b_payload_id,
  output reg  [1:0]    io_axi_b_payload_resp,
  input  wire          io_axi_ar_valid,
  output reg           io_axi_ar_ready,
  input  wire [31:0]   io_axi_ar_payload_addr,
  input  wire [6:0]    io_axi_ar_payload_id,
  input  wire [7:0]    io_axi_ar_payload_len,
  input  wire [2:0]    io_axi_ar_payload_size,
  input  wire [1:0]    io_axi_ar_payload_burst,
  output reg           io_axi_r_valid,
  input  wire          io_axi_r_ready,
  output reg  [31:0]   io_axi_r_payload_data,
  output reg  [6:0]    io_axi_r_payload_id,
  output reg  [1:0]    io_axi_r_payload_resp,
  output reg           io_axi_r_payload_last,
  input  wire [31:0]   io_ram_data_read,
  output wire [31:0]   io_ram_data_write,
  output wire          io_ram_data_writeEnable,
  output wire [19:0]   io_ram_addr,
  output wire [3:0]    io_ram_be_n,
  output wire          io_ram_ce_n,
  output wire          io_ram_oe_n,
  output wire          io_ram_we_n,
  input  wire          clk,
  input  wire          reset
);
  localparam fsm_BOOT = 4'd0;
  localparam fsm_IDLE = 4'd1;
  localparam fsm_VALIDATE = 4'd2;
  localparam fsm_WRITE_DATA_FETCH = 4'd3;
  localparam fsm_WRITE_EXECUTE = 4'd4;
  localparam fsm_WRITE_DEASSERT = 4'd5;
  localparam fsm_WRITE_FINALIZE = 4'd6;
  localparam fsm_WRITE_DATA_ERROR_CONSUME = 4'd7;
  localparam fsm_WRITE_RESPONSE = 4'd8;
  localparam fsm_READ_SETUP = 4'd9;
  localparam fsm_READ_WAIT = 4'd10;
  localparam fsm_READ_RESPONSE = 4'd11;
  localparam fsm_READ_RESPONSE_ERROR = 4'd12;

  wire       [7:0]    _zz_fsm_burst_count_remaining;
  wire       [17:0]   _zz_fsm_current_sram_addr;
  wire       [32:0]   _zz_fsm_current_sram_addr_1;
  wire       [32:0]   _zz_fsm_current_sram_addr_2;
  wire       [7:0]    _zz_fsm_burst_count_remaining_1;
  wire       [17:0]   _zz_fsm_current_sram_addr_3;
  wire       [32:0]   _zz_fsm_current_sram_addr_4;
  wire       [32:0]   _zz_fsm_current_sram_addr_5;
  wire       [19:0]   _zz_fsm_current_sram_addr_6;
  wire       [7:0]    _zz_fsm_current_sram_addr_7;
  wire       [7:0]    _zz_fsm_current_sram_addr_8;
  wire       [19:0]   _zz_fsm_next_sram_addr_prefetch;
  wire       [7:0]    _zz_fsm_next_sram_addr_prefetch_1;
  wire       [7:0]    _zz_fsm_next_sram_addr_prefetch_2;
  wire       [19:0]   _zz_fsm_current_sram_addr_9;
  wire       [7:0]    _zz_fsm_current_sram_addr_10;
  wire       [7:0]    _zz_fsm_current_sram_addr_11;
  wire       [3:0]    sram_be_n_inactive_value;
  (* mark_debug = "TRUE" *) reg        [19:0]   sram_addr_out_reg;
  (* mark_debug = "TRUE" *) reg        [31:0]   sram_data_out_reg;
  (* mark_debug = "TRUE" *) reg        [3:0]    sram_be_n_out_reg;
  (* mark_debug = "TRUE" *) reg                 sram_ce_n_out_reg;
  (* mark_debug = "TRUE" *) reg                 sram_oe_n_out_reg;
  (* mark_debug = "TRUE" *) reg                 sram_we_n_out_reg;
  (* mark_debug = "TRUE" *) reg                 sram_data_writeEnable_out_reg;
  (* mark_debug = "TRUE" *) reg        [31:0]   write_data_buffer;
  (* mark_debug = "TRUE" *) reg        [3:0]    write_strb_buffer;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  (* mark_debug = "TRUE" *) reg        [31:0]   fsm_ar_cmd_reg_addr;
  (* mark_debug = "TRUE" *) reg        [6:0]    fsm_ar_cmd_reg_id;
  (* mark_debug = "TRUE" *) reg        [7:0]    fsm_ar_cmd_reg_len;
  (* mark_debug = "TRUE" *) reg        [2:0]    fsm_ar_cmd_reg_size;
  (* mark_debug = "TRUE" *) reg        [1:0]    fsm_ar_cmd_reg_burst;
  (* mark_debug = "TRUE" *) reg        [31:0]   fsm_aw_cmd_reg_addr;
  (* mark_debug = "TRUE" *) reg        [6:0]    fsm_aw_cmd_reg_id;
  (* mark_debug = "TRUE" *) reg        [7:0]    fsm_aw_cmd_reg_len;
  (* mark_debug = "TRUE" *) reg        [2:0]    fsm_aw_cmd_reg_size;
  (* mark_debug = "TRUE" *) reg        [1:0]    fsm_aw_cmd_reg_burst;
  (* mark_debug = "TRUE" *) reg        [8:0]    fsm_burst_count_remaining;
  (* mark_debug = "TRUE" *) reg        [19:0]   fsm_current_sram_addr;
  (* mark_debug = "TRUE" *) reg        [31:0]   fsm_read_data_buffer;
  reg        [1:0]    fsm_read_wait_counter;
  reg        [1:0]    fsm_write_wait_counter;
  (* MARK_DEBUG = "TRUE" *) reg                 fsm_transaction_error_occurred;
  reg                 fsm_read_priority;
  reg        [19:0]   fsm_next_sram_addr_prefetch;
  reg                 fsm_addr_prefetch_valid;
  (* MARK_DEBUG = "TRUE" *) reg        [3:0]    fsm_stateReg;
  reg        [3:0]    fsm_stateNext;
  wire                when_SRAMController_l293;
  (* mark_debug = "true" *) wire                io_axi_aw_fire;
  (* mark_debug = "true" *) wire                io_axi_ar_fire;
  (* mark_debug = "true" *) wire                io_axi_w_fire;
  wire                when_SRAMController_l454;
  wire                when_SRAMController_l473;
  wire                when_SRAMController_l490;
  wire                when_SRAMController_l523;
  wire                when_SRAMController_l625;
  wire                when_SRAMController_l634;
  wire                when_SRAMController_l664;
  (* mark_debug = "true" *) wire                io_axi_r_fire;
  wire                when_SRAMController_l713;
  wire                fsm_onExit_BOOT;
  wire                fsm_onExit_IDLE;
  wire                fsm_onExit_VALIDATE;
  wire                fsm_onExit_WRITE_DATA_FETCH;
  wire                fsm_onExit_WRITE_EXECUTE;
  wire                fsm_onExit_WRITE_DEASSERT;
  wire                fsm_onExit_WRITE_FINALIZE;
  wire                fsm_onExit_WRITE_DATA_ERROR_CONSUME;
  wire                fsm_onExit_WRITE_RESPONSE;
  wire                fsm_onExit_READ_SETUP;
  wire                fsm_onExit_READ_WAIT;
  wire                fsm_onExit_READ_RESPONSE;
  wire                fsm_onExit_READ_RESPONSE_ERROR;
  wire                fsm_onEntry_BOOT;
  wire                fsm_onEntry_IDLE;
  wire                fsm_onEntry_VALIDATE;
  wire                fsm_onEntry_WRITE_DATA_FETCH;
  wire                fsm_onEntry_WRITE_EXECUTE;
  wire                fsm_onEntry_WRITE_DEASSERT;
  wire                fsm_onEntry_WRITE_FINALIZE;
  wire                fsm_onEntry_WRITE_DATA_ERROR_CONSUME;
  wire                fsm_onEntry_WRITE_RESPONSE;
  wire                fsm_onEntry_READ_SETUP;
  wire                fsm_onEntry_READ_WAIT;
  wire                fsm_onEntry_READ_RESPONSE;
  wire                fsm_onEntry_READ_RESPONSE_ERROR;
  (* mark_debug = "true" *) wire                io_axi_b_fire;
  reg                 sram_ce_n_out_reg_prev;
  reg                 sram_we_n_out_reg_prev;
  wire                when_SRAMController_l749;
  wire                when_SRAMController_l750;
  `ifndef SYNTHESIS
  reg [191:0] fsm_stateReg_string;
  reg [191:0] fsm_stateNext_string;
  `endif


  assign _zz_fsm_burst_count_remaining = (io_axi_aw_payload_len + 8'h01);
  assign _zz_fsm_current_sram_addr = (_zz_fsm_current_sram_addr_1[19 : 0] >>> 2'd2);
  assign _zz_fsm_current_sram_addr_1 = (_zz_fsm_current_sram_addr_2 - 33'h080000000);
  assign _zz_fsm_current_sram_addr_2 = {1'd0, io_axi_aw_payload_addr};
  assign _zz_fsm_burst_count_remaining_1 = (io_axi_ar_payload_len + 8'h01);
  assign _zz_fsm_current_sram_addr_3 = (_zz_fsm_current_sram_addr_4[19 : 0] >>> 2'd2);
  assign _zz_fsm_current_sram_addr_4 = (_zz_fsm_current_sram_addr_5 - 33'h080000000);
  assign _zz_fsm_current_sram_addr_5 = {1'd0, io_axi_ar_payload_addr};
  assign _zz_fsm_current_sram_addr_7 = (_zz_fsm_current_sram_addr_8 / 3'b100);
  assign _zz_fsm_current_sram_addr_6 = {12'd0, _zz_fsm_current_sram_addr_7};
  assign _zz_fsm_current_sram_addr_8 = ({7'd0,1'b1} <<< fsm_aw_cmd_reg_size);
  assign _zz_fsm_next_sram_addr_prefetch_1 = (_zz_fsm_next_sram_addr_prefetch_2 / 3'b100);
  assign _zz_fsm_next_sram_addr_prefetch = {12'd0, _zz_fsm_next_sram_addr_prefetch_1};
  assign _zz_fsm_next_sram_addr_prefetch_2 = ({7'd0,1'b1} <<< fsm_ar_cmd_reg_size);
  assign _zz_fsm_current_sram_addr_10 = (_zz_fsm_current_sram_addr_11 / 3'b100);
  assign _zz_fsm_current_sram_addr_9 = {12'd0, _zz_fsm_current_sram_addr_10};
  assign _zz_fsm_current_sram_addr_11 = ({7'd0,1'b1} <<< fsm_ar_cmd_reg_size);
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_BOOT : fsm_stateReg_string = "BOOT                    ";
      fsm_IDLE : fsm_stateReg_string = "IDLE                    ";
      fsm_VALIDATE : fsm_stateReg_string = "VALIDATE                ";
      fsm_WRITE_DATA_FETCH : fsm_stateReg_string = "WRITE_DATA_FETCH        ";
      fsm_WRITE_EXECUTE : fsm_stateReg_string = "WRITE_EXECUTE           ";
      fsm_WRITE_DEASSERT : fsm_stateReg_string = "WRITE_DEASSERT          ";
      fsm_WRITE_FINALIZE : fsm_stateReg_string = "WRITE_FINALIZE          ";
      fsm_WRITE_DATA_ERROR_CONSUME : fsm_stateReg_string = "WRITE_DATA_ERROR_CONSUME";
      fsm_WRITE_RESPONSE : fsm_stateReg_string = "WRITE_RESPONSE          ";
      fsm_READ_SETUP : fsm_stateReg_string = "READ_SETUP              ";
      fsm_READ_WAIT : fsm_stateReg_string = "READ_WAIT               ";
      fsm_READ_RESPONSE : fsm_stateReg_string = "READ_RESPONSE           ";
      fsm_READ_RESPONSE_ERROR : fsm_stateReg_string = "READ_RESPONSE_ERROR     ";
      default : fsm_stateReg_string = "????????????????????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_BOOT : fsm_stateNext_string = "BOOT                    ";
      fsm_IDLE : fsm_stateNext_string = "IDLE                    ";
      fsm_VALIDATE : fsm_stateNext_string = "VALIDATE                ";
      fsm_WRITE_DATA_FETCH : fsm_stateNext_string = "WRITE_DATA_FETCH        ";
      fsm_WRITE_EXECUTE : fsm_stateNext_string = "WRITE_EXECUTE           ";
      fsm_WRITE_DEASSERT : fsm_stateNext_string = "WRITE_DEASSERT          ";
      fsm_WRITE_FINALIZE : fsm_stateNext_string = "WRITE_FINALIZE          ";
      fsm_WRITE_DATA_ERROR_CONSUME : fsm_stateNext_string = "WRITE_DATA_ERROR_CONSUME";
      fsm_WRITE_RESPONSE : fsm_stateNext_string = "WRITE_RESPONSE          ";
      fsm_READ_SETUP : fsm_stateNext_string = "READ_SETUP              ";
      fsm_READ_WAIT : fsm_stateNext_string = "READ_WAIT               ";
      fsm_READ_RESPONSE : fsm_stateNext_string = "READ_RESPONSE           ";
      fsm_READ_RESPONSE_ERROR : fsm_stateNext_string = "READ_RESPONSE_ERROR     ";
      default : fsm_stateNext_string = "????????????????????????";
    endcase
  end
  `endif

  always @(*) begin
    io_axi_aw_ready = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
        io_axi_aw_ready = 1'b0;
        if(when_SRAMController_l293) begin
          io_axi_aw_ready = (! fsm_read_priority);
        end else begin
          io_axi_aw_ready = io_axi_aw_valid;
        end
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        io_axi_aw_ready = 1'b0;
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_ar_ready = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
        io_axi_ar_ready = 1'b0;
        if(when_SRAMController_l293) begin
          io_axi_ar_ready = fsm_read_priority;
        end else begin
          io_axi_ar_ready = io_axi_ar_valid;
        end
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        io_axi_ar_ready = 1'b0;
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_w_ready = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
        io_axi_w_ready = 1'b0;
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
        io_axi_w_ready = 1'b1;
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        io_axi_w_ready = 1'b1;
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_b_valid = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
        io_axi_b_valid = 1'b1;
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_valid = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_valid = 1'b1;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_b_payload_id = 7'h0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
        io_axi_b_payload_id = fsm_aw_cmd_reg_id;
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_b_payload_resp = 2'b00;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
        io_axi_b_payload_resp = (fsm_transaction_error_occurred ? 2'b10 : 2'b00);
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_payload_id = 7'h0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_payload_id = fsm_ar_cmd_reg_id;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_payload_id = fsm_ar_cmd_reg_id;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_payload_data = 32'h0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_payload_data = fsm_read_data_buffer;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_payload_data = 32'h0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_payload_resp = 2'b00;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_payload_resp = 2'b00;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_payload_resp = 2'b10;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_r_payload_last = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
        io_axi_r_payload_last = when_SRAMController_l664;
      end
      fsm_READ_RESPONSE_ERROR : begin
        io_axi_r_payload_last = when_SRAMController_l713;
      end
      default : begin
      end
    endcase
  end

  assign sram_be_n_inactive_value = 4'b1111;
  assign io_ram_addr = sram_addr_out_reg;
  assign io_ram_ce_n = sram_ce_n_out_reg;
  assign io_ram_oe_n = sram_oe_n_out_reg;
  assign io_ram_we_n = sram_we_n_out_reg;
  assign io_ram_be_n = sram_be_n_out_reg;
  assign io_ram_data_write = sram_data_out_reg;
  assign io_ram_data_writeEnable = sram_data_writeEnable_out_reg;
  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_IDLE : begin
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
      end
      fsm_READ_WAIT : begin
      end
      fsm_READ_RESPONSE : begin
      end
      fsm_READ_RESPONSE_ERROR : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_IDLE : begin
        if(io_axi_aw_fire) begin
          fsm_stateNext = fsm_WRITE_DATA_FETCH;
        end
        if(io_axi_ar_fire) begin
          fsm_stateNext = fsm_READ_SETUP;
        end
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
        if(io_axi_w_fire) begin
          fsm_stateNext = fsm_WRITE_EXECUTE;
        end
      end
      fsm_WRITE_EXECUTE : begin
        if(when_SRAMController_l454) begin
          fsm_stateNext = fsm_WRITE_DEASSERT;
        end
      end
      fsm_WRITE_DEASSERT : begin
        if(when_SRAMController_l473) begin
          fsm_stateNext = fsm_WRITE_FINALIZE;
        end
      end
      fsm_WRITE_FINALIZE : begin
        if(when_SRAMController_l490) begin
          fsm_stateNext = fsm_WRITE_RESPONSE;
        end else begin
          fsm_stateNext = fsm_WRITE_DATA_FETCH;
        end
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        if(io_axi_w_fire) begin
          if(when_SRAMController_l523) begin
            fsm_stateNext = fsm_WRITE_RESPONSE;
          end
        end
      end
      fsm_WRITE_RESPONSE : begin
        if(io_axi_b_ready) begin
          fsm_stateNext = fsm_IDLE;
        end
      end
      fsm_READ_SETUP : begin
        fsm_stateNext = fsm_READ_WAIT;
      end
      fsm_READ_WAIT : begin
        if(when_SRAMController_l634) begin
          fsm_stateNext = fsm_READ_RESPONSE;
        end
      end
      fsm_READ_RESPONSE : begin
        if(io_axi_r_fire) begin
          if(when_SRAMController_l664) begin
            fsm_stateNext = fsm_IDLE;
          end else begin
            fsm_stateNext = fsm_READ_SETUP;
          end
        end
      end
      fsm_READ_RESPONSE_ERROR : begin
        if(io_axi_r_fire) begin
          if(when_SRAMController_l713) begin
            fsm_stateNext = fsm_IDLE;
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_IDLE;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_BOOT;
    end
  end

  assign when_SRAMController_l293 = (io_axi_aw_valid && io_axi_ar_valid);
  assign io_axi_aw_fire = (io_axi_aw_valid && io_axi_aw_ready);
  assign io_axi_ar_fire = (io_axi_ar_valid && io_axi_ar_ready);
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign when_SRAMController_l454 = (fsm_write_wait_counter == 2'b11);
  assign when_SRAMController_l473 = 1'b1;
  assign when_SRAMController_l490 = (fsm_burst_count_remaining == 9'h0);
  assign when_SRAMController_l523 = (fsm_burst_count_remaining == 9'h001);
  assign when_SRAMController_l625 = (((fsm_read_wait_counter == 2'b10) && (9'h001 < fsm_burst_count_remaining)) && (! fsm_addr_prefetch_valid));
  assign when_SRAMController_l634 = (fsm_read_wait_counter == 2'b11);
  assign when_SRAMController_l664 = (fsm_burst_count_remaining == 9'h001);
  assign io_axi_r_fire = (io_axi_r_valid && io_axi_r_ready);
  assign when_SRAMController_l713 = (fsm_burst_count_remaining == 9'h001);
  assign fsm_onExit_BOOT = ((fsm_stateNext != fsm_BOOT) && (fsm_stateReg == fsm_BOOT));
  assign fsm_onExit_IDLE = ((fsm_stateNext != fsm_IDLE) && (fsm_stateReg == fsm_IDLE));
  assign fsm_onExit_VALIDATE = ((fsm_stateNext != fsm_VALIDATE) && (fsm_stateReg == fsm_VALIDATE));
  assign fsm_onExit_WRITE_DATA_FETCH = ((fsm_stateNext != fsm_WRITE_DATA_FETCH) && (fsm_stateReg == fsm_WRITE_DATA_FETCH));
  assign fsm_onExit_WRITE_EXECUTE = ((fsm_stateNext != fsm_WRITE_EXECUTE) && (fsm_stateReg == fsm_WRITE_EXECUTE));
  assign fsm_onExit_WRITE_DEASSERT = ((fsm_stateNext != fsm_WRITE_DEASSERT) && (fsm_stateReg == fsm_WRITE_DEASSERT));
  assign fsm_onExit_WRITE_FINALIZE = ((fsm_stateNext != fsm_WRITE_FINALIZE) && (fsm_stateReg == fsm_WRITE_FINALIZE));
  assign fsm_onExit_WRITE_DATA_ERROR_CONSUME = ((fsm_stateNext != fsm_WRITE_DATA_ERROR_CONSUME) && (fsm_stateReg == fsm_WRITE_DATA_ERROR_CONSUME));
  assign fsm_onExit_WRITE_RESPONSE = ((fsm_stateNext != fsm_WRITE_RESPONSE) && (fsm_stateReg == fsm_WRITE_RESPONSE));
  assign fsm_onExit_READ_SETUP = ((fsm_stateNext != fsm_READ_SETUP) && (fsm_stateReg == fsm_READ_SETUP));
  assign fsm_onExit_READ_WAIT = ((fsm_stateNext != fsm_READ_WAIT) && (fsm_stateReg == fsm_READ_WAIT));
  assign fsm_onExit_READ_RESPONSE = ((fsm_stateNext != fsm_READ_RESPONSE) && (fsm_stateReg == fsm_READ_RESPONSE));
  assign fsm_onExit_READ_RESPONSE_ERROR = ((fsm_stateNext != fsm_READ_RESPONSE_ERROR) && (fsm_stateReg == fsm_READ_RESPONSE_ERROR));
  assign fsm_onEntry_BOOT = ((fsm_stateNext == fsm_BOOT) && (fsm_stateReg != fsm_BOOT));
  assign fsm_onEntry_IDLE = ((fsm_stateNext == fsm_IDLE) && (fsm_stateReg != fsm_IDLE));
  assign fsm_onEntry_VALIDATE = ((fsm_stateNext == fsm_VALIDATE) && (fsm_stateReg != fsm_VALIDATE));
  assign fsm_onEntry_WRITE_DATA_FETCH = ((fsm_stateNext == fsm_WRITE_DATA_FETCH) && (fsm_stateReg != fsm_WRITE_DATA_FETCH));
  assign fsm_onEntry_WRITE_EXECUTE = ((fsm_stateNext == fsm_WRITE_EXECUTE) && (fsm_stateReg != fsm_WRITE_EXECUTE));
  assign fsm_onEntry_WRITE_DEASSERT = ((fsm_stateNext == fsm_WRITE_DEASSERT) && (fsm_stateReg != fsm_WRITE_DEASSERT));
  assign fsm_onEntry_WRITE_FINALIZE = ((fsm_stateNext == fsm_WRITE_FINALIZE) && (fsm_stateReg != fsm_WRITE_FINALIZE));
  assign fsm_onEntry_WRITE_DATA_ERROR_CONSUME = ((fsm_stateNext == fsm_WRITE_DATA_ERROR_CONSUME) && (fsm_stateReg != fsm_WRITE_DATA_ERROR_CONSUME));
  assign fsm_onEntry_WRITE_RESPONSE = ((fsm_stateNext == fsm_WRITE_RESPONSE) && (fsm_stateReg != fsm_WRITE_RESPONSE));
  assign fsm_onEntry_READ_SETUP = ((fsm_stateNext == fsm_READ_SETUP) && (fsm_stateReg != fsm_READ_SETUP));
  assign fsm_onEntry_READ_WAIT = ((fsm_stateNext == fsm_READ_WAIT) && (fsm_stateReg != fsm_READ_WAIT));
  assign fsm_onEntry_READ_RESPONSE = ((fsm_stateNext == fsm_READ_RESPONSE) && (fsm_stateReg != fsm_READ_RESPONSE));
  assign fsm_onEntry_READ_RESPONSE_ERROR = ((fsm_stateNext == fsm_READ_RESPONSE_ERROR) && (fsm_stateReg != fsm_READ_RESPONSE_ERROR));
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  assign when_SRAMController_l749 = ((sram_ce_n_out_reg_prev == 1'b0) && (sram_we_n_out_reg_prev == 1'b0));
  assign when_SRAMController_l750 = ((sram_ce_n_out_reg == 1'b1) && (sram_we_n_out_reg == 1'b1));
  always @(posedge clk) begin
    if(reset) begin
      sram_addr_out_reg <= 20'h0;
      sram_data_out_reg <= 32'h0;
      sram_be_n_out_reg <= sram_be_n_inactive_value;
      sram_ce_n_out_reg <= 1'b1;
      sram_oe_n_out_reg <= 1'b1;
      sram_we_n_out_reg <= 1'b1;
      sram_data_writeEnable_out_reg <= 1'b0;
      fsm_transaction_error_occurred <= 1'b0;
      fsm_read_priority <= 1'b0;
      fsm_addr_prefetch_valid <= 1'b0;
      fsm_stateReg <= fsm_BOOT;
      sram_ce_n_out_reg_prev <= 1'b1;
      sram_we_n_out_reg_prev <= 1'b1;
    end else begin
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_IDLE : begin
          fsm_transaction_error_occurred <= 1'b0;
          fsm_addr_prefetch_valid <= 1'b0;
          if(io_axi_aw_fire) begin
            fsm_read_priority <= (! fsm_read_priority);
            fsm_transaction_error_occurred <= 1'b0;
          end
          if(io_axi_ar_fire) begin
            fsm_read_priority <= (! fsm_read_priority);
            fsm_transaction_error_occurred <= 1'b0;
          end
        end
        fsm_VALIDATE : begin
        end
        fsm_WRITE_DATA_FETCH : begin
        end
        fsm_WRITE_EXECUTE : begin
        end
        fsm_WRITE_DEASSERT : begin
        end
        fsm_WRITE_FINALIZE : begin
        end
        fsm_WRITE_DATA_ERROR_CONSUME : begin
        end
        fsm_WRITE_RESPONSE : begin
        end
        fsm_READ_SETUP : begin
          fsm_addr_prefetch_valid <= 1'b0;
          sram_ce_n_out_reg <= 1'b0;
          sram_oe_n_out_reg <= 1'b0;
          sram_we_n_out_reg <= 1'b1;
          sram_data_writeEnable_out_reg <= 1'b0;
          sram_addr_out_reg <= fsm_current_sram_addr;
          sram_be_n_out_reg <= 4'b0000;
        end
        fsm_READ_WAIT : begin
          if(when_SRAMController_l625) begin
            fsm_addr_prefetch_valid <= 1'b1;
          end
        end
        fsm_READ_RESPONSE : begin
          if(io_axi_r_fire) begin
            if(!when_SRAMController_l664) begin
              if(fsm_addr_prefetch_valid) begin
                fsm_addr_prefetch_valid <= 1'b0;
              end
            end
          end
        end
        fsm_READ_RESPONSE_ERROR : begin
        end
        default : begin
        end
      endcase
      if(fsm_onExit_READ_RESPONSE) begin
        sram_oe_n_out_reg <= 1'b1;
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= sram_be_n_inactive_value;
        sram_addr_out_reg <= 20'h0;
      end
      if(fsm_onEntry_IDLE) begin
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
        sram_oe_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= sram_be_n_inactive_value;
        sram_addr_out_reg <= 20'h0;
      end
      if(fsm_onEntry_WRITE_DATA_FETCH) begin
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
      end
      if(fsm_onEntry_WRITE_EXECUTE) begin
        sram_addr_out_reg <= fsm_current_sram_addr;
        sram_data_out_reg <= io_axi_w_payload_data;
        sram_data_writeEnable_out_reg <= 1'b1;
        sram_be_n_out_reg <= (~ io_axi_w_payload_strb);
        sram_ce_n_out_reg <= 1'b0;
        sram_oe_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b0;
      end
      if(fsm_onEntry_WRITE_DEASSERT) begin
        sram_we_n_out_reg <= 1'b1;
      end
      if(fsm_onEntry_WRITE_FINALIZE) begin
        sram_ce_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
      end
      if(fsm_onEntry_WRITE_DATA_ERROR_CONSUME) begin
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
        sram_oe_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= sram_be_n_inactive_value;
        sram_addr_out_reg <= 20'h0;
      end
      if(fsm_onEntry_WRITE_RESPONSE) begin
        sram_ce_n_out_reg <= 1'b1;
        sram_we_n_out_reg <= 1'b1;
        sram_oe_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= sram_be_n_inactive_value;
        sram_addr_out_reg <= 20'h0;
      end
      if(fsm_onEntry_READ_SETUP) begin
        sram_ce_n_out_reg <= 1'b0;
        sram_oe_n_out_reg <= 1'b0;
        sram_we_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_addr_out_reg <= fsm_current_sram_addr;
        sram_be_n_out_reg <= 4'b0000;
      end
      if(fsm_onEntry_READ_WAIT) begin
        sram_ce_n_out_reg <= 1'b0;
        sram_oe_n_out_reg <= 1'b0;
        sram_we_n_out_reg <= 1'b1;
        sram_data_writeEnable_out_reg <= 1'b0;
        sram_be_n_out_reg <= 4'b0000;
      end
      sram_ce_n_out_reg_prev <= sram_ce_n_out_reg;
      sram_we_n_out_reg_prev <= sram_we_n_out_reg;
      if(when_SRAMController_l749) begin
        if(when_SRAMController_l750) begin
          `ifndef SYNTHESIS
            `ifdef FORMAL
              assert(1'b0); // SRAMController.scala:L751
            `else
              if(!1'b0) begin
                $display("FAILURE This is a bug."); // SRAMController.scala:L751
                $finish;
              end
            `endif
          `endif
        end
      end
    end
  end

  always @(posedge clk) begin
    case(fsm_stateReg)
      fsm_IDLE : begin
        if(io_axi_aw_fire) begin
          fsm_aw_cmd_reg_addr <= io_axi_aw_payload_addr;
          fsm_aw_cmd_reg_id <= io_axi_aw_payload_id;
          fsm_aw_cmd_reg_len <= io_axi_aw_payload_len;
          fsm_aw_cmd_reg_size <= io_axi_aw_payload_size;
          fsm_aw_cmd_reg_burst <= io_axi_aw_payload_burst;
          fsm_burst_count_remaining <= {1'd0, _zz_fsm_burst_count_remaining};
          fsm_current_sram_addr <= {2'd0, _zz_fsm_current_sram_addr};
        end
        if(io_axi_ar_fire) begin
          fsm_ar_cmd_reg_addr <= io_axi_ar_payload_addr;
          fsm_ar_cmd_reg_id <= io_axi_ar_payload_id;
          fsm_ar_cmd_reg_len <= io_axi_ar_payload_len;
          fsm_ar_cmd_reg_size <= io_axi_ar_payload_size;
          fsm_ar_cmd_reg_burst <= io_axi_ar_payload_burst;
          fsm_burst_count_remaining <= {1'd0, _zz_fsm_burst_count_remaining_1};
          fsm_current_sram_addr <= {2'd0, _zz_fsm_current_sram_addr_3};
          fsm_read_wait_counter <= 2'b00;
        end
      end
      fsm_VALIDATE : begin
      end
      fsm_WRITE_DATA_FETCH : begin
      end
      fsm_WRITE_EXECUTE : begin
        if(when_SRAMController_l454) begin
          fsm_burst_count_remaining <= (fsm_burst_count_remaining - 9'h001);
        end else begin
          fsm_write_wait_counter <= (fsm_write_wait_counter + 2'b01);
        end
      end
      fsm_WRITE_DEASSERT : begin
      end
      fsm_WRITE_FINALIZE : begin
        if(!when_SRAMController_l490) begin
          fsm_current_sram_addr <= (fsm_current_sram_addr + _zz_fsm_current_sram_addr_6);
        end
      end
      fsm_WRITE_DATA_ERROR_CONSUME : begin
        if(io_axi_w_fire) begin
          fsm_burst_count_remaining <= (fsm_burst_count_remaining - 9'h001);
        end
      end
      fsm_WRITE_RESPONSE : begin
      end
      fsm_READ_SETUP : begin
        fsm_read_wait_counter <= 2'b00;
      end
      fsm_READ_WAIT : begin
        if(when_SRAMController_l625) begin
          fsm_next_sram_addr_prefetch <= (fsm_current_sram_addr + _zz_fsm_next_sram_addr_prefetch);
        end
        if(when_SRAMController_l634) begin
          fsm_read_data_buffer <= io_ram_data_read;
        end else begin
          fsm_read_wait_counter <= (fsm_read_wait_counter + 2'b01);
        end
      end
      fsm_READ_RESPONSE : begin
        if(io_axi_r_fire) begin
          fsm_burst_count_remaining <= (fsm_burst_count_remaining - 9'h001);
          if(!when_SRAMController_l664) begin
            if(fsm_addr_prefetch_valid) begin
              fsm_current_sram_addr <= fsm_next_sram_addr_prefetch;
            end else begin
              fsm_current_sram_addr <= (fsm_current_sram_addr + _zz_fsm_current_sram_addr_9);
            end
          end
        end
      end
      fsm_READ_RESPONSE_ERROR : begin
        if(io_axi_r_fire) begin
          fsm_burst_count_remaining <= (fsm_burst_count_remaining - 9'h001);
        end
      end
      default : begin
      end
    endcase
    if(fsm_onEntry_WRITE_EXECUTE) begin
      fsm_write_wait_counter <= 2'b00;
    end
  end


endmodule

module IntAlu (
  input  wire          io_iqEntryIn_valid,
  input  wire [3:0]    io_iqEntryIn_payload_robPtr,
  input  wire [5:0]    io_iqEntryIn_payload_physDest_idx,
  input  wire          io_iqEntryIn_payload_physDestIsFpr,
  input  wire          io_iqEntryIn_payload_writesToPhysReg,
  input  wire          io_iqEntryIn_payload_useSrc1,
  input  wire [31:0]   io_iqEntryIn_payload_src1Data,
  input  wire [5:0]    io_iqEntryIn_payload_src1Tag,
  input  wire          io_iqEntryIn_payload_src1Ready,
  input  wire          io_iqEntryIn_payload_src1IsFpr,
  input  wire          io_iqEntryIn_payload_useSrc2,
  input  wire [31:0]   io_iqEntryIn_payload_src2Data,
  input  wire [5:0]    io_iqEntryIn_payload_src2Tag,
  input  wire          io_iqEntryIn_payload_src2Ready,
  input  wire          io_iqEntryIn_payload_src2IsFpr,
  input  wire          io_iqEntryIn_payload_aluCtrl_valid,
  input  wire          io_iqEntryIn_payload_aluCtrl_isSub,
  input  wire          io_iqEntryIn_payload_aluCtrl_isAdd,
  input  wire          io_iqEntryIn_payload_aluCtrl_isSigned,
  input  wire [1:0]    io_iqEntryIn_payload_aluCtrl_logicOp,
  input  wire          io_iqEntryIn_payload_shiftCtrl_valid,
  input  wire          io_iqEntryIn_payload_shiftCtrl_isRight,
  input  wire          io_iqEntryIn_payload_shiftCtrl_isArithmetic,
  input  wire          io_iqEntryIn_payload_shiftCtrl_isRotate,
  input  wire          io_iqEntryIn_payload_shiftCtrl_isDoubleWord,
  input  wire [31:0]   io_iqEntryIn_payload_imm,
  input  wire [2:0]    io_iqEntryIn_payload_immUsage,
  output wire          io_resultOut_valid,
  output reg  [31:0]   io_resultOut_payload_data,
  output reg  [5:0]    io_resultOut_payload_physDest_idx,
  output reg           io_resultOut_payload_writesToPhysReg,
  output reg  [3:0]    io_resultOut_payload_robPtr,
  output reg           io_resultOut_payload_hasException,
  output reg  [0:0]    io_resultOut_payload_exceptionCode
);
  localparam LogicOp_NONE = 2'd0;
  localparam LogicOp_AND_1 = 2'd1;
  localparam LogicOp_OR_1 = 2'd2;
  localparam LogicOp_XOR_1 = 2'd3;
  localparam ImmUsageType_NONE = 3'd0;
  localparam ImmUsageType_SRC_ALU = 3'd1;
  localparam ImmUsageType_SRC_SHIFT_AMT = 3'd2;
  localparam ImmUsageType_SRC_CSR_UIMM = 3'd3;
  localparam ImmUsageType_MEM_OFFSET = 3'd4;
  localparam ImmUsageType_BRANCH_OFFSET = 3'd5;
  localparam ImmUsageType_JUMP_OFFSET = 3'd6;
  localparam IntAluExceptionCode_NONE = 1'd0;
  localparam IntAluExceptionCode_UNDEFINED_ALU_OP = 1'd1;

  wire       [31:0]   _zz_io_resultOut_payload_data_3;
  wire                _zz_io_resultOut_payload_data_4;
  wire       [31:0]   _zz_io_resultOut_payload_data_5;
  wire       [31:0]   _zz_io_resultOut_payload_data_6;
  wire                _zz_io_resultOut_payload_data_7;
  wire       [31:0]   _zz_io_resultOut_payload_data_8;
  wire       [31:0]   _zz_io_resultOut_payload_data_9;
  wire                _zz_io_resultOut_payload_data_10;
  wire       [31:0]   _zz_io_resultOut_payload_data_11;
  wire       [31:0]   _zz_io_resultOut_payload_data_12;
  wire       [31:0]   _zz_io_resultOut_payload_data_13;
  wire       [1:0]    _zz_io_resultOut_payload_data_14;
  wire       [31:0]   _zz_io_resultOut_payload_data_15;
  wire                _zz_io_resultOut_payload_data_16;
  wire       [31:0]   _zz_io_resultOut_payload_data_17;
  wire                _zz_io_resultOut_payload_data_18;
  wire       [31:0]   _zz_io_resultOut_payload_data_19;
  wire       [62:0]   _zz_io_resultOut_payload_data_20;
  wire       [31:0]   _zz_io_resultOut_payload_data_21;
  wire       [31:0]   _zz_io_resultOut_payload_data_22;
  wire       [31:0]   _zz_io_resultOut_payload_data_23;
  wire       [4:0]    _zz_io_resultOut_payload_data;
  wire       [31:0]   _zz_io_resultOut_payload_data_1;
  wire                _zz_io_resultOut_payload_data_2;
  wire       [0:0]    _zz_io_resultOut_payload_exceptionCode;
  `ifndef SYNTHESIS
  reg [39:0] io_iqEntryIn_payload_aluCtrl_logicOp_string;
  reg [103:0] io_iqEntryIn_payload_immUsage_string;
  reg [127:0] io_resultOut_payload_exceptionCode_string;
  reg [127:0] _zz_io_resultOut_payload_exceptionCode_string;
  `endif


  assign _zz_io_resultOut_payload_data_6 = (io_iqEntryIn_payload_src1Data + io_iqEntryIn_payload_src2Data);
  assign _zz_io_resultOut_payload_data_9 = (io_iqEntryIn_payload_src1Data - io_iqEntryIn_payload_src2Data);
  assign _zz_io_resultOut_payload_data_12 = io_iqEntryIn_payload_src1Data;
  assign _zz_io_resultOut_payload_data_13 = io_iqEntryIn_payload_src2Data;
  assign _zz_io_resultOut_payload_data_20 = ({31'd0,io_iqEntryIn_payload_src1Data} <<< _zz_io_resultOut_payload_data);
  assign _zz_io_resultOut_payload_data_19 = _zz_io_resultOut_payload_data_20[31:0];
  assign _zz_io_resultOut_payload_data_21 = (io_iqEntryIn_payload_src1Data >>> _zz_io_resultOut_payload_data);
  assign _zz_io_resultOut_payload_data_22 = ($signed(_zz_io_resultOut_payload_data_23) >>> _zz_io_resultOut_payload_data);
  assign _zz_io_resultOut_payload_data_23 = io_iqEntryIn_payload_src1Data;
  assign _zz_io_resultOut_payload_data_3 = ((((_zz_io_resultOut_payload_data_4 ? _zz_io_resultOut_payload_data_5 : _zz_io_resultOut_payload_data_1) | (_zz_io_resultOut_payload_data_7 ? _zz_io_resultOut_payload_data_8 : _zz_io_resultOut_payload_data_1)) | ((_zz_io_resultOut_payload_data_10 && io_iqEntryIn_payload_aluCtrl_isSigned) ? _zz_io_resultOut_payload_data_11 : _zz_io_resultOut_payload_data_1)) | ((io_iqEntryIn_payload_aluCtrl_valid && (io_iqEntryIn_payload_aluCtrl_logicOp == _zz_io_resultOut_payload_data_14)) ? (io_iqEntryIn_payload_src1Data & io_iqEntryIn_payload_src2Data) : _zz_io_resultOut_payload_data_1));
  assign _zz_io_resultOut_payload_data_15 = ((io_iqEntryIn_payload_aluCtrl_valid && (io_iqEntryIn_payload_aluCtrl_logicOp == LogicOp_OR_1)) ? (io_iqEntryIn_payload_src1Data | io_iqEntryIn_payload_src2Data) : _zz_io_resultOut_payload_data_1);
  assign _zz_io_resultOut_payload_data_16 = (io_iqEntryIn_payload_aluCtrl_valid && (io_iqEntryIn_payload_aluCtrl_logicOp == LogicOp_XOR_1));
  assign _zz_io_resultOut_payload_data_17 = (io_iqEntryIn_payload_src1Data ^ io_iqEntryIn_payload_src2Data);
  assign _zz_io_resultOut_payload_data_18 = (! io_iqEntryIn_payload_shiftCtrl_isRight);
  assign _zz_io_resultOut_payload_data_4 = (io_iqEntryIn_payload_aluCtrl_valid && io_iqEntryIn_payload_aluCtrl_isAdd);
  assign _zz_io_resultOut_payload_data_5 = _zz_io_resultOut_payload_data_6;
  assign _zz_io_resultOut_payload_data_7 = ((io_iqEntryIn_payload_aluCtrl_valid && io_iqEntryIn_payload_aluCtrl_isSub) && (! io_iqEntryIn_payload_aluCtrl_isSigned));
  assign _zz_io_resultOut_payload_data_8 = _zz_io_resultOut_payload_data_9;
  assign _zz_io_resultOut_payload_data_10 = (io_iqEntryIn_payload_aluCtrl_valid && io_iqEntryIn_payload_aluCtrl_isSub);
  assign _zz_io_resultOut_payload_data_11 = (($signed(_zz_io_resultOut_payload_data_12) < $signed(_zz_io_resultOut_payload_data_13)) ? 32'h00000001 : 32'h0);
  assign _zz_io_resultOut_payload_data_14 = LogicOp_AND_1;
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_iqEntryIn_payload_aluCtrl_logicOp)
      LogicOp_NONE : io_iqEntryIn_payload_aluCtrl_logicOp_string = "NONE ";
      LogicOp_AND_1 : io_iqEntryIn_payload_aluCtrl_logicOp_string = "AND_1";
      LogicOp_OR_1 : io_iqEntryIn_payload_aluCtrl_logicOp_string = "OR_1 ";
      LogicOp_XOR_1 : io_iqEntryIn_payload_aluCtrl_logicOp_string = "XOR_1";
      default : io_iqEntryIn_payload_aluCtrl_logicOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_iqEntryIn_payload_immUsage)
      ImmUsageType_NONE : io_iqEntryIn_payload_immUsage_string = "NONE         ";
      ImmUsageType_SRC_ALU : io_iqEntryIn_payload_immUsage_string = "SRC_ALU      ";
      ImmUsageType_SRC_SHIFT_AMT : io_iqEntryIn_payload_immUsage_string = "SRC_SHIFT_AMT";
      ImmUsageType_SRC_CSR_UIMM : io_iqEntryIn_payload_immUsage_string = "SRC_CSR_UIMM ";
      ImmUsageType_MEM_OFFSET : io_iqEntryIn_payload_immUsage_string = "MEM_OFFSET   ";
      ImmUsageType_BRANCH_OFFSET : io_iqEntryIn_payload_immUsage_string = "BRANCH_OFFSET";
      ImmUsageType_JUMP_OFFSET : io_iqEntryIn_payload_immUsage_string = "JUMP_OFFSET  ";
      default : io_iqEntryIn_payload_immUsage_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(io_resultOut_payload_exceptionCode)
      IntAluExceptionCode_NONE : io_resultOut_payload_exceptionCode_string = "NONE            ";
      IntAluExceptionCode_UNDEFINED_ALU_OP : io_resultOut_payload_exceptionCode_string = "UNDEFINED_ALU_OP";
      default : io_resultOut_payload_exceptionCode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_resultOut_payload_exceptionCode)
      IntAluExceptionCode_NONE : _zz_io_resultOut_payload_exceptionCode_string = "NONE            ";
      IntAluExceptionCode_UNDEFINED_ALU_OP : _zz_io_resultOut_payload_exceptionCode_string = "UNDEFINED_ALU_OP";
      default : _zz_io_resultOut_payload_exceptionCode_string = "????????????????";
    endcase
  end
  `endif

  assign io_resultOut_valid = io_iqEntryIn_valid;
  always @(*) begin
    io_resultOut_payload_data = 32'h0;
    if(io_iqEntryIn_valid) begin
      io_resultOut_payload_data = ((! _zz_io_resultOut_payload_data_2) ? _zz_io_resultOut_payload_data_1 : (((((_zz_io_resultOut_payload_data_3 | _zz_io_resultOut_payload_data_15) | (_zz_io_resultOut_payload_data_16 ? _zz_io_resultOut_payload_data_17 : _zz_io_resultOut_payload_data_1)) | ((io_iqEntryIn_payload_shiftCtrl_valid && _zz_io_resultOut_payload_data_18) ? _zz_io_resultOut_payload_data_19 : _zz_io_resultOut_payload_data_1)) | (((io_iqEntryIn_payload_shiftCtrl_valid && io_iqEntryIn_payload_shiftCtrl_isRight) && (! io_iqEntryIn_payload_shiftCtrl_isArithmetic)) ? _zz_io_resultOut_payload_data_21 : _zz_io_resultOut_payload_data_1)) | (((io_iqEntryIn_payload_shiftCtrl_valid && io_iqEntryIn_payload_shiftCtrl_isRight) && io_iqEntryIn_payload_shiftCtrl_isArithmetic) ? _zz_io_resultOut_payload_data_22 : _zz_io_resultOut_payload_data_1)));
    end
  end

  always @(*) begin
    io_resultOut_payload_physDest_idx = 6'h0;
    if(io_iqEntryIn_valid) begin
      io_resultOut_payload_physDest_idx = io_iqEntryIn_payload_physDest_idx;
    end
  end

  always @(*) begin
    io_resultOut_payload_writesToPhysReg = 1'b0;
    if(io_iqEntryIn_valid) begin
      io_resultOut_payload_writesToPhysReg = io_iqEntryIn_payload_writesToPhysReg;
    end
  end

  always @(*) begin
    io_resultOut_payload_robPtr = 4'b0000;
    if(io_iqEntryIn_valid) begin
      io_resultOut_payload_robPtr = io_iqEntryIn_payload_robPtr;
    end
  end

  always @(*) begin
    io_resultOut_payload_hasException = 1'b0;
    if(io_iqEntryIn_valid) begin
      io_resultOut_payload_hasException = (! _zz_io_resultOut_payload_data_2);
    end
  end

  always @(*) begin
    io_resultOut_payload_exceptionCode = IntAluExceptionCode_NONE;
    if(io_iqEntryIn_valid) begin
      io_resultOut_payload_exceptionCode = _zz_io_resultOut_payload_exceptionCode;
    end
  end

  assign _zz_io_resultOut_payload_data = ((io_iqEntryIn_payload_immUsage == ImmUsageType_SRC_SHIFT_AMT) ? io_iqEntryIn_payload_imm[4 : 0] : io_iqEntryIn_payload_src2Data[4 : 0]);
  assign _zz_io_resultOut_payload_data_1 = 32'h0;
  assign _zz_io_resultOut_payload_data_2 = (io_iqEntryIn_payload_aluCtrl_valid || io_iqEntryIn_payload_shiftCtrl_valid);
  assign _zz_io_resultOut_payload_exceptionCode = ((! _zz_io_resultOut_payload_data_2) ? IntAluExceptionCode_UNDEFINED_ALU_OP : IntAluExceptionCode_NONE);

endmodule

//StreamFifoLowLatency_2 replaced by StreamFifoLowLatency

//StreamArbiter_5 replaced by StreamArbiter

//StreamArbiter_4 replaced by StreamArbiter

//StreamFifoLowLatency_1 replaced by StreamFifoLowLatency

//StreamArbiter_3 replaced by StreamArbiter

//StreamArbiter_2 replaced by StreamArbiter

module StreamFifoLowLatency (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [1:0]    io_push_payload,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [1:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire                fifo_io_push_ready;
  wire                fifo_io_pop_valid;
  wire       [1:0]    fifo_io_pop_payload;
  wire       [2:0]    fifo_io_occupancy;
  wire       [2:0]    fifo_io_availability;

  StreamFifo_8 fifo (
    .io_push_valid   (io_push_valid            ), //i
    .io_push_ready   (fifo_io_push_ready       ), //o
    .io_push_payload (io_push_payload[1:0]     ), //i
    .io_pop_valid    (fifo_io_pop_valid        ), //o
    .io_pop_ready    (io_pop_ready             ), //i
    .io_pop_payload  (fifo_io_pop_payload[1:0] ), //o
    .io_flush        (io_flush                 ), //i
    .io_occupancy    (fifo_io_occupancy[2:0]   ), //o
    .io_availability (fifo_io_availability[2:0]), //o
    .clk             (clk                      ), //i
    .reset           (reset                    )  //i
  );
  assign io_push_ready = fifo_io_push_ready;
  assign io_pop_valid = fifo_io_pop_valid;
  assign io_pop_payload = fifo_io_pop_payload;
  assign io_occupancy = fifo_io_occupancy;
  assign io_availability = fifo_io_availability;

endmodule

//StreamArbiter_1 replaced by StreamArbiter

module StreamArbiter (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [31:0]   io_inputs_0_payload_addr,
  input  wire [4:0]    io_inputs_0_payload_id,
  input  wire [7:0]    io_inputs_0_payload_len,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire [1:0]    io_inputs_0_payload_burst,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [31:0]   io_inputs_1_payload_addr,
  input  wire [4:0]    io_inputs_1_payload_id,
  input  wire [7:0]    io_inputs_1_payload_len,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire [1:0]    io_inputs_1_payload_burst,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [31:0]   io_inputs_2_payload_addr,
  input  wire [4:0]    io_inputs_2_payload_id,
  input  wire [7:0]    io_inputs_2_payload_len,
  input  wire [2:0]    io_inputs_2_payload_size,
  input  wire [1:0]    io_inputs_2_payload_burst,
  input  wire          io_inputs_3_valid,
  output wire          io_inputs_3_ready,
  input  wire [31:0]   io_inputs_3_payload_addr,
  input  wire [4:0]    io_inputs_3_payload_id,
  input  wire [7:0]    io_inputs_3_payload_len,
  input  wire [2:0]    io_inputs_3_payload_size,
  input  wire [1:0]    io_inputs_3_payload_burst,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [31:0]   io_output_payload_addr,
  output wire [4:0]    io_output_payload_id,
  output wire [7:0]    io_output_payload_len,
  output wire [2:0]    io_output_payload_size,
  output wire [1:0]    io_output_payload_burst,
  output wire [1:0]    io_chosen,
  output wire [3:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [7:0]    _zz__zz_maskProposal_0_2;
  wire       [7:0]    _zz__zz_maskProposal_0_2_1;
  wire       [3:0]    _zz__zz_maskProposal_0_2_2;
  reg        [31:0]   _zz_io_output_payload_addr_3;
  reg        [4:0]    _zz_io_output_payload_id;
  reg        [7:0]    _zz_io_output_payload_len;
  reg        [2:0]    _zz_io_output_payload_size;
  reg        [1:0]    _zz_io_output_payload_burst;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  wire                maskProposal_3;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  reg                 maskLocked_3;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire                maskRouted_3;
  wire       [3:0]    _zz_maskProposal_0;
  wire       [7:0]    _zz_maskProposal_0_1;
  wire       [7:0]    _zz_maskProposal_0_2;
  wire       [3:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                _zz_io_output_payload_addr;
  wire                _zz_io_output_payload_addr_1;
  wire       [1:0]    _zz_io_output_payload_addr_2;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  wire                _zz_io_chosen_2;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_2,{maskLocked_1,{maskLocked_0,maskLocked_3}}};
  assign _zz__zz_maskProposal_0_2_1 = {4'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(_zz_io_output_payload_addr_2)
      2'b00 : begin
        _zz_io_output_payload_addr_3 = io_inputs_0_payload_addr;
        _zz_io_output_payload_id = io_inputs_0_payload_id;
        _zz_io_output_payload_len = io_inputs_0_payload_len;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_burst = io_inputs_0_payload_burst;
      end
      2'b01 : begin
        _zz_io_output_payload_addr_3 = io_inputs_1_payload_addr;
        _zz_io_output_payload_id = io_inputs_1_payload_id;
        _zz_io_output_payload_len = io_inputs_1_payload_len;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_burst = io_inputs_1_payload_burst;
      end
      2'b10 : begin
        _zz_io_output_payload_addr_3 = io_inputs_2_payload_addr;
        _zz_io_output_payload_id = io_inputs_2_payload_id;
        _zz_io_output_payload_len = io_inputs_2_payload_len;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_burst = io_inputs_2_payload_burst;
      end
      default : begin
        _zz_io_output_payload_addr_3 = io_inputs_3_payload_addr;
        _zz_io_output_payload_id = io_inputs_3_payload_id;
        _zz_io_output_payload_len = io_inputs_3_payload_len;
        _zz_io_output_payload_size = io_inputs_3_payload_size;
        _zz_io_output_payload_burst = io_inputs_3_payload_burst;
      end
    endcase
  end

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign maskRouted_3 = (locked ? maskLocked_3 : maskProposal_3);
  assign _zz_maskProposal_0 = {io_inputs_3_valid,{io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[7 : 4] | _zz_maskProposal_0_2[3 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign maskProposal_3 = _zz_maskProposal_0_3[3];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2)) || (io_inputs_3_valid && maskRouted_3));
  assign _zz_io_output_payload_addr = (maskRouted_1 || maskRouted_3);
  assign _zz_io_output_payload_addr_1 = (maskRouted_2 || maskRouted_3);
  assign _zz_io_output_payload_addr_2 = {_zz_io_output_payload_addr_1,_zz_io_output_payload_addr};
  assign io_output_payload_addr = _zz_io_output_payload_addr_3;
  assign io_output_payload_id = _zz_io_output_payload_id;
  assign io_output_payload_len = _zz_io_output_payload_len;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_burst = _zz_io_output_payload_burst;
  assign io_inputs_0_ready = ((1'b0 || maskRouted_0) && io_output_ready);
  assign io_inputs_1_ready = ((1'b0 || maskRouted_1) && io_output_ready);
  assign io_inputs_2_ready = ((1'b0 || maskRouted_2) && io_output_ready);
  assign io_inputs_3_ready = ((1'b0 || maskRouted_3) && io_output_ready);
  assign io_chosenOH = {maskRouted_3,{maskRouted_2,{maskRouted_1,maskRouted_0}}};
  assign _zz_io_chosen = io_chosenOH[3];
  assign _zz_io_chosen_1 = (io_chosenOH[1] || _zz_io_chosen);
  assign _zz_io_chosen_2 = (io_chosenOH[2] || _zz_io_chosen);
  assign io_chosen = {_zz_io_chosen_2,_zz_io_chosen_1};
  always @(posedge clk) begin
    if(reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b0;
      maskLocked_3 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
        maskLocked_3 <= maskRouted_3;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

//Axi4WriteOnlyErrorSlave_3 replaced by Axi4WriteOnlyErrorSlave

//Axi4ReadOnlyErrorSlave_3 replaced by Axi4ReadOnlyErrorSlave

module Axi4WriteOnlyErrorSlave_2 (
  input  wire          io_axi_aw_valid,
  output wire          io_axi_aw_ready,
  input  wire [31:0]   io_axi_aw_payload_addr,
  input  wire [2:0]    io_axi_aw_payload_id,
  input  wire [7:0]    io_axi_aw_payload_len,
  input  wire [2:0]    io_axi_aw_payload_size,
  input  wire [1:0]    io_axi_aw_payload_burst,
  input  wire [2:0]    io_axi_aw_payload_prot,
  input  wire          io_axi_w_valid,
  output wire          io_axi_w_ready,
  input  wire [31:0]   io_axi_w_payload_data,
  input  wire [3:0]    io_axi_w_payload_strb,
  input  wire          io_axi_w_payload_last,
  output wire          io_axi_b_valid,
  input  wire          io_axi_b_ready,
  output wire [2:0]    io_axi_b_payload_id,
  output wire [1:0]    io_axi_b_payload_resp,
  input  wire          clk,
  input  wire          reset
);

  reg                 consumeData;
  reg                 sendRsp;
  reg        [2:0]    id;
  wire                io_axi_aw_fire;
  wire                io_axi_w_fire;
  wire                when_Axi4ErrorSlave_l24;
  wire                io_axi_b_fire;

  assign io_axi_aw_ready = (! (consumeData || sendRsp));
  assign io_axi_aw_fire = (io_axi_aw_valid && io_axi_aw_ready);
  assign io_axi_w_ready = consumeData;
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign when_Axi4ErrorSlave_l24 = (io_axi_w_fire && io_axi_w_payload_last);
  assign io_axi_b_valid = sendRsp;
  assign io_axi_b_payload_resp = 2'b11;
  assign io_axi_b_payload_id = id;
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  always @(posedge clk) begin
    if(reset) begin
      consumeData <= 1'b0;
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_aw_fire) begin
        consumeData <= 1'b1;
      end
      if(when_Axi4ErrorSlave_l24) begin
        consumeData <= 1'b0;
        sendRsp <= 1'b1;
      end
      if(io_axi_b_fire) begin
        sendRsp <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_axi_aw_fire) begin
      id <= io_axi_aw_payload_id;
    end
  end


endmodule

module Axi4ReadOnlyErrorSlave_2 (
  input  wire          io_axi_ar_valid,
  output wire          io_axi_ar_ready,
  input  wire [31:0]   io_axi_ar_payload_addr,
  input  wire [2:0]    io_axi_ar_payload_id,
  input  wire [7:0]    io_axi_ar_payload_len,
  input  wire [2:0]    io_axi_ar_payload_size,
  input  wire [1:0]    io_axi_ar_payload_burst,
  input  wire [2:0]    io_axi_ar_payload_prot,
  output wire          io_axi_r_valid,
  input  wire          io_axi_r_ready,
  output wire [31:0]   io_axi_r_payload_data,
  output wire [2:0]    io_axi_r_payload_id,
  output wire [1:0]    io_axi_r_payload_resp,
  output wire          io_axi_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  reg                 sendRsp;
  reg        [2:0]    id;
  reg        [7:0]    remaining;
  wire                remainingZero;
  wire                io_axi_ar_fire;

  assign remainingZero = (remaining == 8'h0);
  assign io_axi_ar_ready = (! sendRsp);
  assign io_axi_ar_fire = (io_axi_ar_valid && io_axi_ar_ready);
  assign io_axi_r_valid = sendRsp;
  assign io_axi_r_payload_id = id;
  assign io_axi_r_payload_resp = 2'b11;
  assign io_axi_r_payload_last = remainingZero;
  always @(posedge clk) begin
    if(reset) begin
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_ar_fire) begin
        sendRsp <= 1'b1;
      end
      if(sendRsp) begin
        if(io_axi_r_ready) begin
          if(remainingZero) begin
            sendRsp <= 1'b0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    if(io_axi_ar_fire) begin
      remaining <= io_axi_ar_payload_len;
      id <= io_axi_ar_payload_id;
    end
    if(sendRsp) begin
      if(io_axi_r_ready) begin
        remaining <= (remaining - 8'h01);
      end
    end
  end


endmodule

//Axi4WriteOnlyErrorSlave_1 replaced by Axi4WriteOnlyErrorSlave

//Axi4ReadOnlyErrorSlave_1 replaced by Axi4ReadOnlyErrorSlave

module Axi4WriteOnlyErrorSlave (
  input  wire          io_axi_aw_valid,
  output wire          io_axi_aw_ready,
  input  wire [31:0]   io_axi_aw_payload_addr,
  input  wire [3:0]    io_axi_aw_payload_id,
  input  wire [7:0]    io_axi_aw_payload_len,
  input  wire [2:0]    io_axi_aw_payload_size,
  input  wire [1:0]    io_axi_aw_payload_burst,
  input  wire          io_axi_w_valid,
  output wire          io_axi_w_ready,
  input  wire [31:0]   io_axi_w_payload_data,
  input  wire [3:0]    io_axi_w_payload_strb,
  input  wire          io_axi_w_payload_last,
  output wire          io_axi_b_valid,
  input  wire          io_axi_b_ready,
  output wire [3:0]    io_axi_b_payload_id,
  output wire [1:0]    io_axi_b_payload_resp,
  input  wire          clk,
  input  wire          reset
);

  reg                 consumeData;
  reg                 sendRsp;
  reg        [3:0]    id;
  wire                io_axi_aw_fire;
  wire                io_axi_w_fire;
  wire                when_Axi4ErrorSlave_l24;
  wire                io_axi_b_fire;

  assign io_axi_aw_ready = (! (consumeData || sendRsp));
  assign io_axi_aw_fire = (io_axi_aw_valid && io_axi_aw_ready);
  assign io_axi_w_ready = consumeData;
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign when_Axi4ErrorSlave_l24 = (io_axi_w_fire && io_axi_w_payload_last);
  assign io_axi_b_valid = sendRsp;
  assign io_axi_b_payload_resp = 2'b11;
  assign io_axi_b_payload_id = id;
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  always @(posedge clk) begin
    if(reset) begin
      consumeData <= 1'b0;
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_aw_fire) begin
        consumeData <= 1'b1;
      end
      if(when_Axi4ErrorSlave_l24) begin
        consumeData <= 1'b0;
        sendRsp <= 1'b1;
      end
      if(io_axi_b_fire) begin
        sendRsp <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_axi_aw_fire) begin
      id <= io_axi_aw_payload_id;
    end
  end


endmodule

module Axi4ReadOnlyErrorSlave (
  input  wire          io_axi_ar_valid,
  output wire          io_axi_ar_ready,
  input  wire [31:0]   io_axi_ar_payload_addr,
  input  wire [3:0]    io_axi_ar_payload_id,
  input  wire [7:0]    io_axi_ar_payload_len,
  input  wire [2:0]    io_axi_ar_payload_size,
  input  wire [1:0]    io_axi_ar_payload_burst,
  output wire          io_axi_r_valid,
  input  wire          io_axi_r_ready,
  output wire [31:0]   io_axi_r_payload_data,
  output wire [3:0]    io_axi_r_payload_id,
  output wire [1:0]    io_axi_r_payload_resp,
  output wire          io_axi_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  reg                 sendRsp;
  reg        [3:0]    id;
  reg        [7:0]    remaining;
  wire                remainingZero;
  wire                io_axi_ar_fire;

  assign remainingZero = (remaining == 8'h0);
  assign io_axi_ar_ready = (! sendRsp);
  assign io_axi_ar_fire = (io_axi_ar_valid && io_axi_ar_ready);
  assign io_axi_r_valid = sendRsp;
  assign io_axi_r_payload_id = id;
  assign io_axi_r_payload_resp = 2'b11;
  assign io_axi_r_payload_last = remainingZero;
  always @(posedge clk) begin
    if(reset) begin
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_ar_fire) begin
        sendRsp <= 1'b1;
      end
      if(sendRsp) begin
        if(io_axi_r_ready) begin
          if(remainingZero) begin
            sendRsp <= 1'b0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    if(io_axi_ar_fire) begin
      remaining <= io_axi_ar_payload_len;
      id <= io_axi_ar_payload_id;
    end
    if(sendRsp) begin
      if(io_axi_r_ready) begin
        remaining <= (remaining - 8'h01);
      end
    end
  end


endmodule

//StreamFifo_7 replaced by StreamFifo_3

//StreamFork_1 replaced by StreamFork

//StreamFifo_6 replaced by StreamFifo_2

//StreamFifo_5 replaced by StreamFifo_1

//StreamFifo_4 replaced by StreamFifo

module StreamFifo_3 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [3:0]    io_push_payload_id,
  input  wire [1:0]    io_push_payload_resp,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [3:0]    io_pop_payload_id,
  output wire [1:0]    io_pop_payload_resp,
  input  wire          io_flush,
  output wire [1:0]    io_occupancy,
  output wire [1:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [5:0]    logic_ram_spinal_port1;
  wire       [5:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [1:0]    logic_ptr_push;
  reg        [1:0]    logic_ptr_pop;
  wire       [1:0]    logic_ptr_occupancy;
  wire       [1:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1455;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [0:0]    logic_push_onRam_write_payload_address;
  wire       [3:0]    logic_push_onRam_write_payload_data_id;
  wire       [1:0]    logic_push_onRam_write_payload_data_resp;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [0:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [0:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [0:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l477;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [0:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [3:0]    logic_pop_sync_readPort_rsp_id;
  wire       [1:0]    logic_pop_sync_readPort_rsp_resp;
  wire       [5:0]    _zz_logic_pop_sync_readPort_rsp_id;
  wire                logic_pop_addressGen_toFlowFire_valid;
  wire       [0:0]    logic_pop_addressGen_toFlowFire_payload;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_id;
  wire       [1:0]    logic_pop_sync_readArbitation_translated_payload_resp;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [1:0]    logic_pop_sync_popReg;
  (* ram_style = "block" *) reg [5:0] logic_ram [0:1];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_resp,logic_push_onRam_write_payload_data_id};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1455 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 2'b10) == 2'b00);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[0:0];
  assign logic_push_onRam_write_payload_data_id = io_push_payload_id;
  assign logic_push_onRam_write_payload_data_resp = io_push_payload_resp;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[0:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l477) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_id = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_id = _zz_logic_pop_sync_readPort_rsp_id[3 : 0];
  assign logic_pop_sync_readPort_rsp_resp = _zz_logic_pop_sync_readPort_rsp_id[5 : 4];
  assign logic_pop_addressGen_toFlowFire_valid = logic_pop_addressGen_fire;
  assign logic_pop_addressGen_toFlowFire_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_toFlowFire_valid;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_toFlowFire_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_id = logic_pop_sync_readPort_rsp_id;
  assign logic_pop_sync_readArbitation_translated_payload_resp = logic_pop_sync_readPort_rsp_resp;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_id = logic_pop_sync_readArbitation_translated_payload_id;
  assign io_pop_payload_resp = logic_pop_sync_readArbitation_translated_payload_resp;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (2'b10 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 2'b00;
      logic_ptr_pop <= 2'b00;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 2'b00;
    end else begin
      if(when_Stream_l1455) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 2'b01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 2'b01);
      end
      if(io_flush) begin
        logic_ptr_push <= 2'b00;
        logic_ptr_pop <= 2'b00;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 2'b00;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module StreamFork (
  input  wire          io_input_valid,
  output reg           io_input_ready,
  input  wire [31:0]   io_input_payload_address,
  input  wire [31:0]   io_input_payload_data,
  input  wire [3:0]    io_input_payload_byteEnables,
  input  wire [3:0]    io_input_payload_id,
  input  wire          io_input_payload_last,
  output wire          io_outputs_0_valid,
  input  wire          io_outputs_0_ready,
  output wire [31:0]   io_outputs_0_payload_address,
  output wire [31:0]   io_outputs_0_payload_data,
  output wire [3:0]    io_outputs_0_payload_byteEnables,
  output wire [3:0]    io_outputs_0_payload_id,
  output wire          io_outputs_0_payload_last,
  output wire          io_outputs_1_valid,
  input  wire          io_outputs_1_ready,
  output wire [31:0]   io_outputs_1_payload_address,
  output wire [31:0]   io_outputs_1_payload_data,
  output wire [3:0]    io_outputs_1_payload_byteEnables,
  output wire [3:0]    io_outputs_1_payload_id,
  output wire          io_outputs_1_payload_last,
  input  wire          clk,
  input  wire          reset
);

  reg                 logic_linkEnable_0;
  reg                 logic_linkEnable_1;
  wire                when_Stream_l1253;
  wire                when_Stream_l1253_1;
  wire                io_outputs_0_fire;
  wire                io_outputs_1_fire;

  always @(*) begin
    io_input_ready = 1'b1;
    if(when_Stream_l1253) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l1253_1) begin
      io_input_ready = 1'b0;
    end
  end

  assign when_Stream_l1253 = ((! io_outputs_0_ready) && logic_linkEnable_0);
  assign when_Stream_l1253_1 = ((! io_outputs_1_ready) && logic_linkEnable_1);
  assign io_outputs_0_valid = (io_input_valid && logic_linkEnable_0);
  assign io_outputs_0_payload_address = io_input_payload_address;
  assign io_outputs_0_payload_data = io_input_payload_data;
  assign io_outputs_0_payload_byteEnables = io_input_payload_byteEnables;
  assign io_outputs_0_payload_id = io_input_payload_id;
  assign io_outputs_0_payload_last = io_input_payload_last;
  assign io_outputs_0_fire = (io_outputs_0_valid && io_outputs_0_ready);
  assign io_outputs_1_valid = (io_input_valid && logic_linkEnable_1);
  assign io_outputs_1_payload_address = io_input_payload_address;
  assign io_outputs_1_payload_data = io_input_payload_data;
  assign io_outputs_1_payload_byteEnables = io_input_payload_byteEnables;
  assign io_outputs_1_payload_id = io_input_payload_id;
  assign io_outputs_1_payload_last = io_input_payload_last;
  assign io_outputs_1_fire = (io_outputs_1_valid && io_outputs_1_ready);
  always @(posedge clk) begin
    if(reset) begin
      logic_linkEnable_0 <= 1'b1;
      logic_linkEnable_1 <= 1'b1;
    end else begin
      if(io_outputs_0_fire) begin
        logic_linkEnable_0 <= 1'b0;
      end
      if(io_outputs_1_fire) begin
        logic_linkEnable_1 <= 1'b0;
      end
      if(io_input_ready) begin
        logic_linkEnable_0 <= 1'b1;
        logic_linkEnable_1 <= 1'b1;
      end
    end
  end


endmodule

module StreamFifo_2 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_address,
  input  wire [31:0]   io_push_payload_data,
  input  wire [3:0]    io_push_payload_byteEnables,
  input  wire [3:0]    io_push_payload_id,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_address,
  output wire [31:0]   io_pop_payload_data,
  output wire [3:0]    io_pop_payload_byteEnables,
  output wire [3:0]    io_pop_payload_id,
  output wire          io_pop_payload_last,
  input  wire          io_flush,
  output wire [1:0]    io_occupancy,
  output wire [1:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [72:0]   logic_ram_spinal_port1;
  wire       [72:0]   _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [1:0]    logic_ptr_push;
  reg        [1:0]    logic_ptr_pop;
  wire       [1:0]    logic_ptr_occupancy;
  wire       [1:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1455;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [0:0]    logic_push_onRam_write_payload_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_data;
  wire       [3:0]    logic_push_onRam_write_payload_data_byteEnables;
  wire       [3:0]    logic_push_onRam_write_payload_data_id;
  wire                logic_push_onRam_write_payload_data_last;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [0:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [0:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [0:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l477;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [0:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [31:0]   logic_pop_sync_readPort_rsp_address;
  wire       [31:0]   logic_pop_sync_readPort_rsp_data;
  wire       [3:0]    logic_pop_sync_readPort_rsp_byteEnables;
  wire       [3:0]    logic_pop_sync_readPort_rsp_id;
  wire                logic_pop_sync_readPort_rsp_last;
  wire       [72:0]   _zz_logic_pop_sync_readPort_rsp_address;
  wire                logic_pop_addressGen_toFlowFire_valid;
  wire       [0:0]    logic_pop_addressGen_toFlowFire_payload;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_address;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_data;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_byteEnables;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_id;
  wire                logic_pop_sync_readArbitation_translated_payload_last;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [1:0]    logic_pop_sync_popReg;
  (* ram_style = "block" *) reg [72:0] logic_ram [0:1];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_last,{logic_push_onRam_write_payload_data_id,{logic_push_onRam_write_payload_data_byteEnables,{logic_push_onRam_write_payload_data_data,logic_push_onRam_write_payload_data_address}}}};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1455 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 2'b10) == 2'b00);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[0:0];
  assign logic_push_onRam_write_payload_data_address = io_push_payload_address;
  assign logic_push_onRam_write_payload_data_data = io_push_payload_data;
  assign logic_push_onRam_write_payload_data_byteEnables = io_push_payload_byteEnables;
  assign logic_push_onRam_write_payload_data_id = io_push_payload_id;
  assign logic_push_onRam_write_payload_data_last = io_push_payload_last;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[0:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l477) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_address = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_address = _zz_logic_pop_sync_readPort_rsp_address[31 : 0];
  assign logic_pop_sync_readPort_rsp_data = _zz_logic_pop_sync_readPort_rsp_address[63 : 32];
  assign logic_pop_sync_readPort_rsp_byteEnables = _zz_logic_pop_sync_readPort_rsp_address[67 : 64];
  assign logic_pop_sync_readPort_rsp_id = _zz_logic_pop_sync_readPort_rsp_address[71 : 68];
  assign logic_pop_sync_readPort_rsp_last = _zz_logic_pop_sync_readPort_rsp_address[72];
  assign logic_pop_addressGen_toFlowFire_valid = logic_pop_addressGen_fire;
  assign logic_pop_addressGen_toFlowFire_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_toFlowFire_valid;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_toFlowFire_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_address = logic_pop_sync_readPort_rsp_address;
  assign logic_pop_sync_readArbitation_translated_payload_data = logic_pop_sync_readPort_rsp_data;
  assign logic_pop_sync_readArbitation_translated_payload_byteEnables = logic_pop_sync_readPort_rsp_byteEnables;
  assign logic_pop_sync_readArbitation_translated_payload_id = logic_pop_sync_readPort_rsp_id;
  assign logic_pop_sync_readArbitation_translated_payload_last = logic_pop_sync_readPort_rsp_last;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_address = logic_pop_sync_readArbitation_translated_payload_address;
  assign io_pop_payload_data = logic_pop_sync_readArbitation_translated_payload_data;
  assign io_pop_payload_byteEnables = logic_pop_sync_readArbitation_translated_payload_byteEnables;
  assign io_pop_payload_id = logic_pop_sync_readArbitation_translated_payload_id;
  assign io_pop_payload_last = logic_pop_sync_readArbitation_translated_payload_last;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (2'b10 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 2'b00;
      logic_ptr_pop <= 2'b00;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 2'b00;
    end else begin
      if(when_Stream_l1455) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 2'b01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 2'b01);
      end
      if(io_flush) begin
        logic_ptr_push <= 2'b00;
        logic_ptr_pop <= 2'b00;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 2'b00;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module StreamFifo_1 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_data,
  input  wire [3:0]    io_push_payload_id,
  input  wire [1:0]    io_push_payload_resp,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_data,
  output wire [3:0]    io_pop_payload_id,
  output wire [1:0]    io_pop_payload_resp,
  output wire          io_pop_payload_last,
  input  wire          io_flush,
  output wire [1:0]    io_occupancy,
  output wire [1:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [38:0]   logic_ram_spinal_port1;
  wire       [38:0]   _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [1:0]    logic_ptr_push;
  reg        [1:0]    logic_ptr_pop;
  wire       [1:0]    logic_ptr_occupancy;
  wire       [1:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1455;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [0:0]    logic_push_onRam_write_payload_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_data;
  wire       [3:0]    logic_push_onRam_write_payload_data_id;
  wire       [1:0]    logic_push_onRam_write_payload_data_resp;
  wire                logic_push_onRam_write_payload_data_last;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [0:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [0:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [0:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l477;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [0:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [31:0]   logic_pop_sync_readPort_rsp_data;
  wire       [3:0]    logic_pop_sync_readPort_rsp_id;
  wire       [1:0]    logic_pop_sync_readPort_rsp_resp;
  wire                logic_pop_sync_readPort_rsp_last;
  wire       [38:0]   _zz_logic_pop_sync_readPort_rsp_data;
  wire                logic_pop_addressGen_toFlowFire_valid;
  wire       [0:0]    logic_pop_addressGen_toFlowFire_payload;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_data;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_id;
  wire       [1:0]    logic_pop_sync_readArbitation_translated_payload_resp;
  wire                logic_pop_sync_readArbitation_translated_payload_last;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [1:0]    logic_pop_sync_popReg;
  (* ram_style = "block" *) reg [38:0] logic_ram [0:1];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_last,{logic_push_onRam_write_payload_data_resp,{logic_push_onRam_write_payload_data_id,logic_push_onRam_write_payload_data_data}}};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1455 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 2'b10) == 2'b00);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[0:0];
  assign logic_push_onRam_write_payload_data_data = io_push_payload_data;
  assign logic_push_onRam_write_payload_data_id = io_push_payload_id;
  assign logic_push_onRam_write_payload_data_resp = io_push_payload_resp;
  assign logic_push_onRam_write_payload_data_last = io_push_payload_last;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[0:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l477) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_data = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_data = _zz_logic_pop_sync_readPort_rsp_data[31 : 0];
  assign logic_pop_sync_readPort_rsp_id = _zz_logic_pop_sync_readPort_rsp_data[35 : 32];
  assign logic_pop_sync_readPort_rsp_resp = _zz_logic_pop_sync_readPort_rsp_data[37 : 36];
  assign logic_pop_sync_readPort_rsp_last = _zz_logic_pop_sync_readPort_rsp_data[38];
  assign logic_pop_addressGen_toFlowFire_valid = logic_pop_addressGen_fire;
  assign logic_pop_addressGen_toFlowFire_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_toFlowFire_valid;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_toFlowFire_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_data = logic_pop_sync_readPort_rsp_data;
  assign logic_pop_sync_readArbitation_translated_payload_id = logic_pop_sync_readPort_rsp_id;
  assign logic_pop_sync_readArbitation_translated_payload_resp = logic_pop_sync_readPort_rsp_resp;
  assign logic_pop_sync_readArbitation_translated_payload_last = logic_pop_sync_readPort_rsp_last;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = logic_pop_sync_readArbitation_translated_payload_data;
  assign io_pop_payload_id = logic_pop_sync_readArbitation_translated_payload_id;
  assign io_pop_payload_resp = logic_pop_sync_readArbitation_translated_payload_resp;
  assign io_pop_payload_last = logic_pop_sync_readArbitation_translated_payload_last;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (2'b10 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 2'b00;
      logic_ptr_pop <= 2'b00;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 2'b00;
    end else begin
      if(when_Stream_l1455) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 2'b01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 2'b01);
      end
      if(io_flush) begin
        logic_ptr_push <= 2'b00;
        logic_ptr_pop <= 2'b00;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 2'b00;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_address,
  input  wire [3:0]    io_push_payload_id,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_address,
  output wire [3:0]    io_pop_payload_id,
  input  wire          io_flush,
  output wire [1:0]    io_occupancy,
  output wire [1:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [35:0]   logic_ram_spinal_port1;
  wire       [35:0]   _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [1:0]    logic_ptr_push;
  reg        [1:0]    logic_ptr_pop;
  wire       [1:0]    logic_ptr_occupancy;
  wire       [1:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1455;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [0:0]    logic_push_onRam_write_payload_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_address;
  wire       [3:0]    logic_push_onRam_write_payload_data_id;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [0:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [0:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [0:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l477;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [0:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [31:0]   logic_pop_sync_readPort_rsp_address;
  wire       [3:0]    logic_pop_sync_readPort_rsp_id;
  wire       [35:0]   _zz_logic_pop_sync_readPort_rsp_address;
  wire                logic_pop_addressGen_toFlowFire_valid;
  wire       [0:0]    logic_pop_addressGen_toFlowFire_payload;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_address;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_id;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [1:0]    logic_pop_sync_popReg;
  (* ram_style = "block" *) reg [35:0] logic_ram [0:1];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_id,logic_push_onRam_write_payload_data_address};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1455 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 2'b10) == 2'b00);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[0:0];
  assign logic_push_onRam_write_payload_data_address = io_push_payload_address;
  assign logic_push_onRam_write_payload_data_id = io_push_payload_id;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[0:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l477) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l477 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_address = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_address = _zz_logic_pop_sync_readPort_rsp_address[31 : 0];
  assign logic_pop_sync_readPort_rsp_id = _zz_logic_pop_sync_readPort_rsp_address[35 : 32];
  assign logic_pop_addressGen_toFlowFire_valid = logic_pop_addressGen_fire;
  assign logic_pop_addressGen_toFlowFire_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_toFlowFire_valid;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_toFlowFire_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_address = logic_pop_sync_readPort_rsp_address;
  assign logic_pop_sync_readArbitation_translated_payload_id = logic_pop_sync_readPort_rsp_id;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_address = logic_pop_sync_readArbitation_translated_payload_address;
  assign io_pop_payload_id = logic_pop_sync_readArbitation_translated_payload_id;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (2'b10 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 2'b00;
      logic_ptr_pop <= 2'b00;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 2'b00;
    end else begin
      if(when_Stream_l1455) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 2'b01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 2'b01);
      end
      if(io_flush) begin
        logic_ptr_push <= 2'b00;
        logic_ptr_pop <= 2'b00;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 2'b00;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

//StreamFifo_10 replaced by StreamFifo_8

//StreamFifo_9 replaced by StreamFifo_8

module StreamFifo_8 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [1:0]    io_push_payload,
  output reg           io_pop_valid,
  input  wire          io_pop_ready,
  output reg  [1:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire       [1:0]    logic_ram_spinal_port1;
  wire       [1:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  reg                 logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1455;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [1:0]    logic_push_onRam_write_payload_address;
  wire       [1:0]    logic_push_onRam_write_payload_data;
  wire                logic_pop_addressGen_valid;
  wire                logic_pop_addressGen_ready;
  wire       [1:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire       [1:0]    logic_pop_async_readed;
  wire                logic_pop_addressGen_translated_valid;
  wire                logic_pop_addressGen_translated_ready;
  wire       [1:0]    logic_pop_addressGen_translated_payload;
  (* ram_style = "distributed" *) reg [1:0] logic_ram [0:3];

  assign _zz_logic_ram_port = logic_push_onRam_write_payload_data;
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  assign logic_ram_spinal_port1 = logic_ram[logic_pop_addressGen_payload];
  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1455 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 3'b100) == 3'b000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  always @(*) begin
    logic_ptr_doPush = io_push_fire;
    if(logic_ptr_empty) begin
      if(io_pop_ready) begin
        logic_ptr_doPush = 1'b0;
      end
    end
  end

  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[1:0];
  assign logic_push_onRam_write_payload_data = io_push_payload;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[1:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  assign logic_pop_async_readed = logic_ram_spinal_port1;
  assign logic_pop_addressGen_translated_valid = logic_pop_addressGen_valid;
  assign logic_pop_addressGen_ready = logic_pop_addressGen_translated_ready;
  assign logic_pop_addressGen_translated_payload = logic_pop_async_readed;
  always @(*) begin
    io_pop_valid = logic_pop_addressGen_translated_valid;
    if(logic_ptr_empty) begin
      io_pop_valid = io_push_valid;
    end
  end

  assign logic_pop_addressGen_translated_ready = io_pop_ready;
  always @(*) begin
    io_pop_payload = logic_pop_addressGen_translated_payload;
    if(logic_ptr_empty) begin
      io_pop_payload = io_push_payload;
    end
  end

  assign logic_ptr_popOnIo = logic_ptr_pop;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b100 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
    end else begin
      if(when_Stream_l1455) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
    end
  end


endmodule
